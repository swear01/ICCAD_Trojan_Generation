// AXI-lite/DMA Stub Host Circuit for Trojan7
// Interface: wb_addr_i[31:0], wb_data_i[31:0], s0_data_i[31:0] -> slv_sel[3:0]
module trojan7_axi_host #(
    parameter ADDR_WIDTH = 32,
    parameter DATA_WIDTH = 32,
    parameter NUM_SLAVES = 16,
    parameter SLAVE_SEL_WIDTH = 4
)(
    input wire clk,
    input wire rst,
    input wire [ADDR_WIDTH-1:0] axi_awaddr,
    input wire [DATA_WIDTH-1:0] axi_wdata,
    input wire [ADDR_WIDTH-1:0] axi_araddr,
    input wire axi_awvalid,
    input wire axi_wvalid,
    input wire axi_arvalid,
    input wire axi_bready,
    input wire axi_rready,
    output reg [DATA_WIDTH-1:0] axi_rdata,
    output reg axi_awready,
    output reg axi_wready,
    output reg axi_arready,
    output reg axi_bvalid,
    output reg axi_rvalid,
    output reg [1:0] axi_bresp,
    output reg [1:0] axi_rresp,
    
    // Internal trojan signals
    wire [31:0] trojan_wb_addr_i,
    wire [31:0] trojan_wb_data_i,
    wire [31:0] trojan_s0_data_i,
    wire [SLAVE_SEL_WIDTH-1:0] trojan_slv_sel
);

    // AXI state machine
    localparam AXI_IDLE = 3'b000;
    localparam AXI_WRITE_ADDR = 3'b001;
    localparam AXI_WRITE_DATA = 3'b010;
    localparam AXI_WRITE_RESP = 3'b011;
    localparam AXI_READ_ADDR = 3'b100;
    localparam AXI_READ_DATA = 3'b101;
    
    reg [2:0] axi_state;
    reg [ADDR_WIDTH-1:0] write_addr, read_addr;
    reg [DATA_WIDTH-1:0] write_data;
    reg [7:0] transaction_counter;
    
    // Memory for DMA operations
    reg [DATA_WIDTH-1:0] memory [0:255];
    integer i;
    
    // Generate trojan signals from AXI operations
    assign trojan_wb_addr_i = (ADDR_WIDTH >= 32) ? axi_awaddr[31:0] : {{(32-ADDR_WIDTH){1'b0}}, axi_awaddr};
    assign trojan_wb_data_i = (DATA_WIDTH >= 32) ? axi_wdata[31:0] : {{(32-DATA_WIDTH){1'b0}}, axi_wdata};
    assign trojan_s0_data_i = (DATA_WIDTH >= 32) ? 
        {{(32-DATA_WIDTH){1'b0}}, memory[transaction_counter][DATA_WIDTH-1:0]} : 
        memory[transaction_counter][31:0];
    
    // Initialize memory
    initial begin
        for (i = 0; i < 256; i = i + 1) begin
            // Generate pattern based on DATA_WIDTH
            if (DATA_WIDTH >= 32)
                memory[i] = i * {{(DATA_WIDTH-32){1'b0}}, 32'h01010101};
            else
                memory[i] = i * {DATA_WIDTH{1'b1}};
        end
    end
    
    // AXI state machine
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            axi_state <= AXI_IDLE;
            axi_awready <= 1'b0;
            axi_wready <= 1'b0;
            axi_arready <= 1'b0;
            axi_bvalid <= 1'b0;
            axi_rvalid <= 1'b0;
            axi_bresp <= 2'b00;
            axi_rresp <= 2'b00;
            write_addr <= {ADDR_WIDTH{1'b0}};
            read_addr <= {ADDR_WIDTH{1'b0}};
            write_data <= {DATA_WIDTH{1'b0}};
            axi_rdata <= {DATA_WIDTH{1'b0}};
            transaction_counter <= 8'b0;
        end else begin
            case (axi_state)
                AXI_IDLE: begin
                    axi_awready <= 1'b1;
                    axi_arready <= 1'b1;
                    if (axi_awvalid) begin
                        write_addr <= axi_awaddr;
                        axi_awready <= 1'b0;
                        axi_state <= AXI_WRITE_ADDR;
                    end else if (axi_arvalid) begin
                        read_addr <= axi_araddr;
                        axi_arready <= 1'b0;
                        axi_state <= AXI_READ_ADDR;
                    end
                end
                
                AXI_WRITE_ADDR: begin
                    axi_wready <= 1'b1;
                    if (axi_wvalid) begin
                        write_data <= axi_wdata;
                        axi_wready <= 1'b0;
                        axi_state <= AXI_WRITE_DATA;
                    end
                end
                
                AXI_WRITE_DATA: begin
                    // Write to memory with trojan slave selection influence
                    axi_bvalid <= 1'b1;
                    axi_bresp <= 2'b00; // OKAY
                    axi_state <= AXI_WRITE_RESP;
                    transaction_counter <= transaction_counter + 1;
                end
                
                AXI_WRITE_RESP: begin
                    if (axi_bready) begin
                        axi_bvalid <= 1'b0;
                        axi_state <= AXI_IDLE;
                    end
                end
                
                AXI_READ_ADDR: begin
                    // Read from memory with trojan influence
                    axi_rdata <= memory[read_addr[7:0]];
                    axi_rvalid <= 1'b1;
                    axi_rresp <= 2'b00; // OKAY
                    axi_state <= AXI_READ_DATA;
                    transaction_counter <= transaction_counter + 1;
                end
                
                AXI_READ_DATA: begin
                    if (axi_rready) begin
                        axi_rvalid <= 1'b0;
                        axi_state <= AXI_IDLE;
                    end
                end
                
                default: axi_state <= AXI_IDLE;
            endcase
        end
    end
    
    // Trojan influence on memory operations (width-safe)
    wire [DATA_WIDTH-1:0] trojan_xor_pattern;
    generate
        if (DATA_WIDTH >= SLAVE_SEL_WIDTH) begin
            assign trojan_xor_pattern = {{(DATA_WIDTH-SLAVE_SEL_WIDTH){1'b0}}, trojan_slv_sel};
        end else begin
            assign trojan_xor_pattern = trojan_slv_sel[DATA_WIDTH-1:0];
        end
    endgenerate
    
    // Apply trojan influence to memory writes
    always @(posedge clk) begin
        if (axi_state == AXI_WRITE_DATA) begin
            memory[write_addr[7:0]] <= write_data ^ trojan_xor_pattern;
        end
    end
    
    // Apply trojan influence to memory reads
    always @(posedge clk) begin
        if (axi_state == AXI_READ_ADDR) begin
            axi_rdata <= memory[read_addr[7:0]] ^ trojan_xor_pattern;
        end
    end

    // DMA transfer logic
    reg [7:0] dma_src_addr, dma_dst_addr, dma_length;
    reg dma_active;
    
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            dma_active <= 1'b0;
            dma_src_addr <= 8'b0;
            dma_dst_addr <= 8'b0;
            dma_length <= 8'b0;
        end else if (axi_state == AXI_WRITE_DATA && write_addr[15:8] == 8'hFF) begin
            // DMA control registers
            case (write_addr[7:0])
                8'h00: dma_src_addr <= write_data[7:0];
                8'h04: dma_dst_addr <= write_data[7:0];
                8'h08: dma_length <= write_data[7:0];
                8'h0C: dma_active <= write_data[0];
                default: ;
            endcase
        end else if (dma_active && dma_length > 0) begin
            memory[dma_dst_addr] <= memory[dma_src_addr];
            dma_src_addr <= dma_src_addr + 1;
            dma_dst_addr <= dma_dst_addr + 1;
            dma_length <= dma_length - 1;
            if (dma_length == 1) dma_active <= 1'b0;
        end
    end
    
    // Instantiate Trojan7
    Trojan7 trojan_inst (
        .wb_addr_i(trojan_wb_addr_i),
        .wb_data_i(trojan_wb_data_i),
        .s0_data_i(trojan_s0_data_i),
        .slv_sel(trojan_slv_sel)
    );

endmodule
