module trojan0_pwm_host_0002(clk, rst, duty_cycle, period, pwm_enable, pwm_out, period_complete);
  wire _000_;
  wire [2:0] _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  input clk;
  wire clk;
  input [7:0] duty_cycle;
  wire [7:0] duty_cycle;
  input [7:0] period;
  wire [7:0] period;
  output period_complete;
  wire period_complete;
  wire [2:0] prescaler_counter;
  wire [7:0] pwm_counter;
  input pwm_enable;
  wire pwm_enable;
  output pwm_out;
  wire pwm_out;
  wire pwm_tick;
  input rst;
  wire rst;
    not _130_(_004_, rst);
    not _131_(_094_, pwm_tick);
    and _132_(_095_, _094_, pwm_counter[0]);
    not _133_(_096_, pwm_counter[0]);
    xor _134_(_097_, period[0], pwm_counter[0]);
    xor _135_(_098_, period[1], pwm_counter[1]);
    or _136_(_099_, _098_, _097_);
    xor _137_(_100_, period[2], pwm_counter[2]);
    xor _138_(_101_, period[3], pwm_counter[3]);
    or _139_(_102_, _101_, _100_);
    or _140_(_103_, _102_, _099_);
    xor _141_(_104_, period[4], pwm_counter[4]);
    xor _142_(_105_, period[5], pwm_counter[5]);
    or _143_(_106_, _105_, _104_);
    xor _144_(_107_, period[6], pwm_counter[6]);
    xor _145_(_108_, period[7], pwm_counter[7]);
    or _146_(_109_, _108_, _107_);
    or _147_(_110_, _109_, _106_);
    or _148_(_111_, _110_, _103_);
    and _149_(_112_, _111_, _096_);
    and _150_(_113_, _112_, pwm_tick);
    or _151_(_018_, _113_, _095_);
    and _152_(_114_, pwm_counter[1], _094_);
    xor _153_(_115_, pwm_counter[1], pwm_counter[0]);
    and _154_(_116_, _115_, _111_);
    and _155_(_117_, _116_, pwm_tick);
    or _156_(_019_, _117_, _114_);
    and _157_(_118_, pwm_counter[2], _094_);
    and _158_(_119_, pwm_counter[1], pwm_counter[0]);
    xor _159_(_120_, _119_, pwm_counter[2]);
    and _160_(_121_, _120_, _111_);
    and _161_(_122_, _121_, pwm_tick);
    or _162_(_020_, _122_, _118_);
    and _163_(_123_, pwm_counter[3], _094_);
    and _164_(_124_, _119_, pwm_counter[2]);
    xor _165_(_125_, _124_, pwm_counter[3]);
    and _166_(_126_, _125_, _111_);
    and _167_(_127_, _126_, pwm_tick);
    or _168_(_021_, _127_, _123_);
    and _169_(_128_, pwm_counter[4], _094_);
    and _170_(_129_, pwm_counter[3], pwm_counter[2]);
    and _171_(_026_, _129_, _119_);
    xor _172_(_027_, _026_, pwm_counter[4]);
    and _173_(_028_, _027_, _111_);
    and _174_(_029_, _028_, pwm_tick);
    or _175_(_022_, _029_, _128_);
    and _176_(_030_, pwm_counter[5], _094_);
    and _177_(_031_, _026_, pwm_counter[4]);
    xor _178_(_032_, _031_, pwm_counter[5]);
    and _179_(_033_, _032_, _111_);
    and _180_(_034_, _033_, pwm_tick);
    or _181_(_023_, _034_, _030_);
    and _182_(_035_, pwm_counter[6], _094_);
    and _183_(_036_, pwm_counter[5], pwm_counter[4]);
    and _184_(_037_, _036_, _026_);
    xor _185_(_038_, _037_, pwm_counter[6]);
    and _186_(_039_, _038_, _111_);
    and _187_(_040_, _039_, pwm_tick);
    or _188_(_024_, _040_, _035_);
    and _189_(_041_, pwm_counter[7], _094_);
    and _190_(_042_, _037_, pwm_counter[6]);
    xor _191_(_043_, _042_, pwm_counter[7]);
    and _192_(_044_, _043_, _111_);
    and _193_(_045_, _044_, pwm_tick);
    or _194_(_025_, _045_, _041_);
    xnor _195_(_046_, duty_cycle[7], pwm_counter[7]);
    xnor _196_(_047_, duty_cycle[6], pwm_counter[6]);
    and _197_(_048_, _047_, _046_);
    xnor _198_(_049_, duty_cycle[5], pwm_counter[5]);
    xnor _199_(_050_, duty_cycle[4], pwm_counter[4]);
    and _200_(_051_, _050_, _049_);
    and _201_(_052_, _051_, _048_);
    xnor _202_(_053_, duty_cycle[3], pwm_counter[3]);
    xnor _203_(_054_, duty_cycle[2], pwm_counter[2]);
    and _204_(_055_, _054_, _053_);
    xnor _205_(_056_, duty_cycle[1], pwm_counter[1]);
    xnor _206_(_057_, duty_cycle[0], pwm_counter[0]);
    and _207_(_058_, _057_, _056_);
    and _208_(_059_, _058_, _055_);
    and _209_(_060_, _059_, _052_);
    not _210_(_061_, pwm_counter[7]);
    and _211_(_062_, duty_cycle[7], _061_);
    not _212_(_063_, pwm_counter[6]);
    and _213_(_064_, duty_cycle[6], _063_);
    and _214_(_065_, _064_, _046_);
    or _215_(_066_, _065_, _062_);
    not _216_(_067_, pwm_counter[5]);
    and _217_(_068_, duty_cycle[5], _067_);
    not _218_(_069_, pwm_counter[4]);
    and _219_(_070_, duty_cycle[4], _069_);
    and _220_(_071_, _070_, _049_);
    or _221_(_072_, _071_, _068_);
    and _222_(_073_, _072_, _048_);
    or _223_(_074_, _073_, _066_);
    not _224_(_075_, pwm_counter[3]);
    and _225_(_076_, duty_cycle[3], _075_);
    not _226_(_077_, pwm_counter[2]);
    and _227_(_078_, duty_cycle[2], _077_);
    and _228_(_079_, _078_, _053_);
    or _229_(_080_, _079_, _076_);
    not _230_(_081_, pwm_counter[1]);
    and _231_(_082_, duty_cycle[1], _081_);
    or _232_(_083_, duty_cycle[0], _096_);
    and _233_(_084_, _083_, _056_);
    or _234_(_085_, _084_, _082_);
    and _235_(_086_, _085_, _055_);
    or _236_(_087_, _086_, _080_);
    and _237_(_088_, _087_, _052_);
    or _238_(_089_, _088_, _074_);
    or _239_(_090_, _089_, _060_);
    and _240_(_002_, _090_, pwm_enable);
    nor _241_(_000_, _111_, _094_);
    and _242_(_091_, prescaler_counter[0], prescaler_counter[1]);
    and _243_(_092_, _091_, prescaler_counter[2]);
    and _244_(_003_, _092_, pwm_enable);
    nor _245_(_001_[0], _092_, prescaler_counter[0]);
    xnor _246_(_093_, prescaler_counter[0], prescaler_counter[1]);
    nor _247_(_001_[1], _093_, _092_);
    xor _248_(_001_[2], _091_, prescaler_counter[2]);
    not _249_(_005_, rst);
    not _250_(_006_, rst);
    not _251_(_007_, rst);
    not _252_(_008_, rst);
    not _253_(_009_, rst);
    not _254_(_010_, rst);
    not _255_(_011_, rst);
    not _256_(_012_, rst);
    not _257_(_013_, rst);
    not _258_(_014_, rst);
    not _259_(_015_, rst);
    not _260_(_016_, rst);
    not _261_(_017_, rst);
    dff _262_(.RN(_004_), .SN(1'b1), .CK(clk), .D(_002_), .Q(pwm_out));
    dff _263_(.RN(_005_), .SN(1'b1), .CK(clk), .D(_000_), .Q(period_complete));
    dff _264_(.RN(_006_), .SN(1'b1), .CK(clk), .D(_001_[0]), .Q(prescaler_counter[0]));
    dff _265_(.RN(_007_), .SN(1'b1), .CK(clk), .D(_001_[1]), .Q(prescaler_counter[1]));
    dff _266_(.RN(_008_), .SN(1'b1), .CK(clk), .D(_001_[2]), .Q(prescaler_counter[2]));
    dff _267_(.RN(_009_), .SN(1'b1), .CK(clk), .D(_003_), .Q(pwm_tick));
    dff _268_(.RN(_010_), .SN(1'b1), .CK(clk), .D(_018_), .Q(pwm_counter[0]));
    dff _269_(.RN(_011_), .SN(1'b1), .CK(clk), .D(_019_), .Q(pwm_counter[1]));
    dff _270_(.RN(_012_), .SN(1'b1), .CK(clk), .D(_020_), .Q(pwm_counter[2]));
    dff _271_(.RN(_013_), .SN(1'b1), .CK(clk), .D(_021_), .Q(pwm_counter[3]));
    dff _272_(.RN(_014_), .SN(1'b1), .CK(clk), .D(_022_), .Q(pwm_counter[4]));
    dff _273_(.RN(_015_), .SN(1'b1), .CK(clk), .D(_023_), .Q(pwm_counter[5]));
    dff _274_(.RN(_016_), .SN(1'b1), .CK(clk), .D(_024_), .Q(pwm_counter[6]));
    dff _275_(.RN(_017_), .SN(1'b1), .CK(clk), .D(_025_), .Q(pwm_counter[7]));
endmodule