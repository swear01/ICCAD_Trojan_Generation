module trojan0_cache_host_0002(clk, rst, addr_tag, addr_index, write_data, cache_read, cache_write, read_data, cache_hit, cache_ready);
  wire _0000_;
  wire _0001_;
  wire _0002_;
  wire _0003_;
  wire _0004_;
  wire _0005_;
  wire _0006_;
  wire _0007_;
  wire _0008_;
  wire _0009_;
  wire _0010_;
  wire _0011_;
  wire _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  wire _0514_;
  wire _0515_;
  wire _0516_;
  wire _0517_;
  wire _0518_;
  wire _0519_;
  wire _0520_;
  wire _0521_;
  wire _0522_;
  wire _0523_;
  wire _0524_;
  wire _0525_;
  wire _0526_;
  wire _0527_;
  wire _0528_;
  wire _0529_;
  wire _0530_;
  wire _0531_;
  wire _0532_;
  wire _0533_;
  wire _0534_;
  wire _0535_;
  wire _0536_;
  wire _0537_;
  wire _0538_;
  wire _0539_;
  wire _0540_;
  wire _0541_;
  wire _0542_;
  wire _0543_;
  wire _0544_;
  wire _0545_;
  wire _0546_;
  wire _0547_;
  wire _0548_;
  wire _0549_;
  wire _0550_;
  wire _0551_;
  wire _0552_;
  wire _0553_;
  wire _0554_;
  wire _0555_;
  wire _0556_;
  wire _0557_;
  wire _0558_;
  wire _0559_;
  wire _0560_;
  wire _0561_;
  wire _0562_;
  wire _0563_;
  wire _0564_;
  wire _0565_;
  wire _0566_;
  wire _0567_;
  wire _0568_;
  wire _0569_;
  wire _0570_;
  wire _0571_;
  wire _0572_;
  wire _0573_;
  wire _0574_;
  wire _0575_;
  wire _0576_;
  wire _0577_;
  wire _0578_;
  wire _0579_;
  wire _0580_;
  wire _0581_;
  wire _0582_;
  wire _0583_;
  wire _0584_;
  wire _0585_;
  wire _0586_;
  wire _0587_;
  wire _0588_;
  wire _0589_;
  wire _0590_;
  wire _0591_;
  wire _0592_;
  wire _0593_;
  wire _0594_;
  wire _0595_;
  wire _0596_;
  wire _0597_;
  wire _0598_;
  wire _0599_;
  wire _0600_;
  wire _0601_;
  wire _0602_;
  wire _0603_;
  wire _0604_;
  wire _0605_;
  wire _0606_;
  wire _0607_;
  wire _0608_;
  wire _0609_;
  wire _0610_;
  wire _0611_;
  wire _0612_;
  wire _0613_;
  wire _0614_;
  wire _0615_;
  wire _0616_;
  wire _0617_;
  wire _0618_;
  wire _0619_;
  wire _0620_;
  wire _0621_;
  wire _0622_;
  wire _0623_;
  wire _0624_;
  wire _0625_;
  wire _0626_;
  wire _0627_;
  wire _0628_;
  wire _0629_;
  wire _0630_;
  wire _0631_;
  wire _0632_;
  wire _0633_;
  wire _0634_;
  wire _0635_;
  wire _0636_;
  wire _0637_;
  wire _0638_;
  wire _0639_;
  wire _0640_;
  wire _0641_;
  wire _0642_;
  wire _0643_;
  wire _0644_;
  wire _0645_;
  wire _0646_;
  wire _0647_;
  wire _0648_;
  wire _0649_;
  wire _0650_;
  wire _0651_;
  wire _0652_;
  wire _0653_;
  wire _0654_;
  wire _0655_;
  wire _0656_;
  wire _0657_;
  wire _0658_;
  wire _0659_;
  wire _0660_;
  wire _0661_;
  wire _0662_;
  wire _0663_;
  wire _0664_;
  wire _0665_;
  wire _0666_;
  wire _0667_;
  wire _0668_;
  wire _0669_;
  wire _0670_;
  wire _0671_;
  wire _0672_;
  wire _0673_;
  wire _0674_;
  wire _0675_;
  wire _0676_;
  wire _0677_;
  wire _0678_;
  wire _0679_;
  wire _0680_;
  wire _0681_;
  wire _0682_;
  wire _0683_;
  wire _0684_;
  wire _0685_;
  wire _0686_;
  wire _0687_;
  wire _0688_;
  wire _0689_;
  wire _0690_;
  wire _0691_;
  wire _0692_;
  wire _0693_;
  wire _0694_;
  wire _0695_;
  wire _0696_;
  wire _0697_;
  wire _0698_;
  wire _0699_;
  wire _0700_;
  wire _0701_;
  wire _0702_;
  wire _0703_;
  wire _0704_;
  wire _0705_;
  wire _0706_;
  wire _0707_;
  wire _0708_;
  wire _0709_;
  wire _0710_;
  wire _0711_;
  wire _0712_;
  wire _0713_;
  wire _0714_;
  wire _0715_;
  wire _0716_;
  wire _0717_;
  wire _0718_;
  wire _0719_;
  wire _0720_;
  wire _0721_;
  wire _0722_;
  wire _0723_;
  wire _0724_;
  wire _0725_;
  wire _0726_;
  wire _0727_;
  wire _0728_;
  wire _0729_;
  wire _0730_;
  wire _0731_;
  wire _0732_;
  wire _0733_;
  wire _0734_;
  wire _0735_;
  wire _0736_;
  wire _0737_;
  wire _0738_;
  wire _0739_;
  wire _0740_;
  wire _0741_;
  wire _0742_;
  wire _0743_;
  wire _0744_;
  wire _0745_;
  wire _0746_;
  wire _0747_;
  wire _0748_;
  wire _0749_;
  wire _0750_;
  wire _0751_;
  wire _0752_;
  wire _0753_;
  wire _0754_;
  wire _0755_;
  wire _0756_;
  wire _0757_;
  wire _0758_;
  wire _0759_;
  wire _0760_;
  wire _0761_;
  wire _0762_;
  wire _0763_;
  wire _0764_;
  wire _0765_;
  wire _0766_;
  wire _0767_;
  wire _0768_;
  wire _0769_;
  wire _0770_;
  wire _0771_;
  wire _0772_;
  wire _0773_;
  wire _0774_;
  wire _0775_;
  wire _0776_;
  wire _0777_;
  wire _0778_;
  wire _0779_;
  wire _0780_;
  wire _0781_;
  wire _0782_;
  wire _0783_;
  wire _0784_;
  wire _0785_;
  wire _0786_;
  wire _0787_;
  wire _0788_;
  wire _0789_;
  wire _0790_;
  wire _0791_;
  wire _0792_;
  wire _0793_;
  wire _0794_;
  wire _0795_;
  wire _0796_;
  wire _0797_;
  wire _0798_;
  wire _0799_;
  wire _0800_;
  wire _0801_;
  wire _0802_;
  wire _0803_;
  wire _0804_;
  wire _0805_;
  wire _0806_;
  wire _0807_;
  wire _0808_;
  wire _0809_;
  wire _0810_;
  wire _0811_;
  wire _0812_;
  wire _0813_;
  wire _0814_;
  wire _0815_;
  wire _0816_;
  wire _0817_;
  wire _0818_;
  wire _0819_;
  wire _0820_;
  wire _0821_;
  wire _0822_;
  wire _0823_;
  wire _0824_;
  wire _0825_;
  wire _0826_;
  wire _0827_;
  wire _0828_;
  wire _0829_;
  wire _0830_;
  wire _0831_;
  wire _0832_;
  wire _0833_;
  wire _0834_;
  wire _0835_;
  wire _0836_;
  wire _0837_;
  wire _0838_;
  wire _0839_;
  wire _0840_;
  wire _0841_;
  wire _0842_;
  wire _0843_;
  wire _0844_;
  wire _0845_;
  wire _0846_;
  wire _0847_;
  wire _0848_;
  wire _0849_;
  wire _0850_;
  wire _0851_;
  wire _0852_;
  wire _0853_;
  wire _0854_;
  wire _0855_;
  wire _0856_;
  wire _0857_;
  wire _0858_;
  wire _0859_;
  wire _0860_;
  wire _0861_;
  wire _0862_;
  wire _0863_;
  wire _0864_;
  wire _0865_;
  wire _0866_;
  wire _0867_;
  wire _0868_;
  wire _0869_;
  wire _0870_;
  wire _0871_;
  wire _0872_;
  wire _0873_;
  wire _0874_;
  wire _0875_;
  wire _0876_;
  wire _0877_;
  wire _0878_;
  wire _0879_;
  wire _0880_;
  wire _0881_;
  wire _0882_;
  wire _0883_;
  wire _0884_;
  wire _0885_;
  wire _0886_;
  wire _0887_;
  wire _0888_;
  wire _0889_;
  wire _0890_;
  wire _0891_;
  wire _0892_;
  wire _0893_;
  wire _0894_;
  wire _0895_;
  wire _0896_;
  wire _0897_;
  wire _0898_;
  wire _0899_;
  wire _0900_;
  wire _0901_;
  wire _0902_;
  wire _0903_;
  wire _0904_;
  wire _0905_;
  wire _0906_;
  wire _0907_;
  wire _0908_;
  wire _0909_;
  wire _0910_;
  wire _0911_;
  wire _0912_;
  wire _0913_;
  wire _0914_;
  wire _0915_;
  wire _0916_;
  wire _0917_;
  wire _0918_;
  wire _0919_;
  wire _0920_;
  wire _0921_;
  wire _0922_;
  wire _0923_;
  wire _0924_;
  wire _0925_;
  wire _0926_;
  wire _0927_;
  wire _0928_;
  wire _0929_;
  wire _0930_;
  wire _0931_;
  wire _0932_;
  wire _0933_;
  wire _0934_;
  wire _0935_;
  wire _0936_;
  wire _0937_;
  wire _0938_;
  wire _0939_;
  wire _0940_;
  wire _0941_;
  wire _0942_;
  wire _0943_;
  wire _0944_;
  wire _0945_;
  wire _0946_;
  wire _0947_;
  wire _0948_;
  wire _0949_;
  wire _0950_;
  wire _0951_;
  wire _0952_;
  wire _0953_;
  wire _0954_;
  wire _0955_;
  wire _0956_;
  wire _0957_;
  wire _0958_;
  wire _0959_;
  wire _0960_;
  wire _0961_;
  wire _0962_;
  wire _0963_;
  wire _0964_;
  wire _0965_;
  wire _0966_;
  wire _0967_;
  wire _0968_;
  wire _0969_;
  wire _0970_;
  wire _0971_;
  wire _0972_;
  wire _0973_;
  wire _0974_;
  wire _0975_;
  wire _0976_;
  wire _0977_;
  wire _0978_;
  wire _0979_;
  wire _0980_;
  wire _0981_;
  wire _0982_;
  wire _0983_;
  wire _0984_;
  wire _0985_;
  wire _0986_;
  wire _0987_;
  wire _0988_;
  wire _0989_;
  wire _0990_;
  wire _0991_;
  wire _0992_;
  wire _0993_;
  wire _0994_;
  wire _0995_;
  wire _0996_;
  wire _0997_;
  wire _0998_;
  wire _0999_;
  wire _1000_;
  wire _1001_;
  wire _1002_;
  wire _1003_;
  wire _1004_;
  wire _1005_;
  wire _1006_;
  wire _1007_;
  wire _1008_;
  wire _1009_;
  wire _1010_;
  wire _1011_;
  wire _1012_;
  wire _1013_;
  wire _1014_;
  wire _1015_;
  wire _1016_;
  wire _1017_;
  wire _1018_;
  wire _1019_;
  wire _1020_;
  wire _1021_;
  wire _1022_;
  wire _1023_;
  wire _1024_;
  wire _1025_;
  wire _1026_;
  wire _1027_;
  wire _1028_;
  wire _1029_;
  wire _1030_;
  wire _1031_;
  wire _1032_;
  wire _1033_;
  wire _1034_;
  wire _1035_;
  wire _1036_;
  wire _1037_;
  wire _1038_;
  wire _1039_;
  wire _1040_;
  wire _1041_;
  wire _1042_;
  wire _1043_;
  wire _1044_;
  wire _1045_;
  wire _1046_;
  wire _1047_;
  wire _1048_;
  wire _1049_;
  wire _1050_;
  wire _1051_;
  wire _1052_;
  wire _1053_;
  wire _1054_;
  wire _1055_;
  wire _1056_;
  wire _1057_;
  wire _1058_;
  wire _1059_;
  wire _1060_;
  wire _1061_;
  wire _1062_;
  wire _1063_;
  wire _1064_;
  wire _1065_;
  wire _1066_;
  wire _1067_;
  wire _1068_;
  wire _1069_;
  wire _1070_;
  wire _1071_;
  wire _1072_;
  wire _1073_;
  wire _1074_;
  wire _1075_;
  wire _1076_;
  wire _1077_;
  wire _1078_;
  wire _1079_;
  wire _1080_;
  wire _1081_;
  wire _1082_;
  wire _1083_;
  wire _1084_;
  wire _1085_;
  wire _1086_;
  wire _1087_;
  wire _1088_;
  wire _1089_;
  wire _1090_;
  wire _1091_;
  wire _1092_;
  wire _1093_;
  wire _1094_;
  wire _1095_;
  wire _1096_;
  wire _1097_;
  wire _1098_;
  wire _1099_;
  wire _1100_;
  wire _1101_;
  wire _1102_;
  wire _1103_;
  wire _1104_;
  wire _1105_;
  wire _1106_;
  wire _1107_;
  wire _1108_;
  wire _1109_;
  wire _1110_;
  wire _1111_;
  wire _1112_;
  wire _1113_;
  wire _1114_;
  wire _1115_;
  wire _1116_;
  wire _1117_;
  wire _1118_;
  wire _1119_;
  wire _1120_;
  wire _1121_;
  wire _1122_;
  wire _1123_;
  wire _1124_;
  wire _1125_;
  wire _1126_;
  wire _1127_;
  wire _1128_;
  wire _1129_;
  wire _1130_;
  wire _1131_;
  wire _1132_;
  wire _1133_;
  wire _1134_;
  wire _1135_;
  wire _1136_;
  wire _1137_;
  wire _1138_;
  wire _1139_;
  wire _1140_;
  wire _1141_;
  wire _1142_;
  wire _1143_;
  wire _1144_;
  wire _1145_;
  wire _1146_;
  wire _1147_;
  wire _1148_;
  wire _1149_;
  wire _1150_;
  wire _1151_;
  wire _1152_;
  wire _1153_;
  wire _1154_;
  wire _1155_;
  wire _1156_;
  wire _1157_;
  wire _1158_;
  wire _1159_;
  wire _1160_;
  wire _1161_;
  wire _1162_;
  wire _1163_;
  wire _1164_;
  wire _1165_;
  wire _1166_;
  wire _1167_;
  wire _1168_;
  wire _1169_;
  wire _1170_;
  wire _1171_;
  wire _1172_;
  wire _1173_;
  wire _1174_;
  wire _1175_;
  wire _1176_;
  wire _1177_;
  wire _1178_;
  wire _1179_;
  wire _1180_;
  wire _1181_;
  wire _1182_;
  wire _1183_;
  wire _1184_;
  wire _1185_;
  wire _1186_;
  wire _1187_;
  wire _1188_;
  wire _1189_;
  wire _1190_;
  wire _1191_;
  wire _1192_;
  wire _1193_;
  wire _1194_;
  wire _1195_;
  wire _1196_;
  wire _1197_;
  wire _1198_;
  wire _1199_;
  wire _1200_;
  wire _1201_;
  wire _1202_;
  wire _1203_;
  wire _1204_;
  wire _1205_;
  wire _1206_;
  wire _1207_;
  wire _1208_;
  wire _1209_;
  wire _1210_;
  wire _1211_;
  wire _1212_;
  wire _1213_;
  wire _1214_;
  wire _1215_;
  wire _1216_;
  wire _1217_;
  wire _1218_;
  wire _1219_;
  wire _1220_;
  wire _1221_;
  wire _1222_;
  wire _1223_;
  wire _1224_;
  wire _1225_;
  wire _1226_;
  wire _1227_;
  wire _1228_;
  wire _1229_;
  wire _1230_;
  wire _1231_;
  wire _1232_;
  wire _1233_;
  wire _1234_;
  wire _1235_;
  wire _1236_;
  wire _1237_;
  wire _1238_;
  wire _1239_;
  wire _1240_;
  wire _1241_;
  wire _1242_;
  wire _1243_;
  wire _1244_;
  wire _1245_;
  wire _1246_;
  wire _1247_;
  wire _1248_;
  wire _1249_;
  wire _1250_;
  wire _1251_;
  wire _1252_;
  wire _1253_;
  wire _1254_;
  wire _1255_;
  wire _1256_;
  wire _1257_;
  wire _1258_;
  wire _1259_;
  wire _1260_;
  wire _1261_;
  wire _1262_;
  wire _1263_;
  wire _1264_;
  wire _1265_;
  wire _1266_;
  wire _1267_;
  wire _1268_;
  wire _1269_;
  wire _1270_;
  wire _1271_;
  wire _1272_;
  wire _1273_;
  wire _1274_;
  wire _1275_;
  wire _1276_;
  wire _1277_;
  wire _1278_;
  wire _1279_;
  wire _1280_;
  wire _1281_;
  wire _1282_;
  wire _1283_;
  wire _1284_;
  wire _1285_;
  wire _1286_;
  wire _1287_;
  wire _1288_;
  wire _1289_;
  wire _1290_;
  wire _1291_;
  wire _1292_;
  wire _1293_;
  wire _1294_;
  wire _1295_;
  wire _1296_;
  wire _1297_;
  wire _1298_;
  wire _1299_;
  wire _1300_;
  wire _1301_;
  wire _1302_;
  wire _1303_;
  wire _1304_;
  wire _1305_;
  wire _1306_;
  wire _1307_;
  wire _1308_;
  wire _1309_;
  wire _1310_;
  wire _1311_;
  wire _1312_;
  wire _1313_;
  wire _1314_;
  wire _1315_;
  wire _1316_;
  wire _1317_;
  wire _1318_;
  wire _1319_;
  wire _1320_;
  wire _1321_;
  wire _1322_;
  wire _1323_;
  wire [2:0] access_index;
  input [5:0] addr_index;
  wire [5:0] addr_index;
  input [3:0] addr_tag;
  wire [3:0] addr_tag;
  wire [15:0] \cache_data[0] ;
  wire [15:0] \cache_data[1] ;
  wire [15:0] \cache_data[2] ;
  wire [15:0] \cache_data[3] ;
  wire [15:0] \cache_data[4] ;
  wire [15:0] \cache_data[5] ;
  wire [15:0] \cache_data[6] ;
  wire [15:0] \cache_data[7] ;
  output cache_hit;
  wire cache_hit;
  input cache_read;
  wire cache_read;
  output cache_ready;
  wire cache_ready;
  wire [2:0] cache_state;
  wire [3:0] \cache_tags[0] ;
  wire [3:0] \cache_tags[1] ;
  wire [3:0] \cache_tags[2] ;
  wire [3:0] \cache_tags[3] ;
  wire [3:0] \cache_tags[4] ;
  wire [3:0] \cache_tags[5] ;
  wire [3:0] \cache_tags[6] ;
  wire [3:0] \cache_tags[7] ;
  input cache_write;
  wire cache_write;
  input clk;
  wire clk;
  output [15:0] read_data;
  wire [15:0] read_data;
  input rst;
  wire rst;
  wire [7:0] valid_bits;
  input [15:0] write_data;
  wire [15:0] write_data;
    not _1324_(_0000_, rst);
    not _1325_(_1044_, cache_state[2]);
    not _1326_(_1045_, cache_state[1]);
    and _1327_(_1046_, _1045_, cache_state[0]);
    and _1328_(_1047_, _1046_, _1044_);
    and _1329_(_1048_, _1047_, cache_write);
    not _1330_(_1049_, access_index[0]);
    and _1331_(_1050_, access_index[1], _1049_);
    and _1332_(_1051_, _1050_, access_index[2]);
    and _1333_(_1052_, _1051_, _1048_);
    not _1334_(_1053_, _1052_);
    and _1335_(_1054_, _1053_, \cache_tags[6][0]);
    and _1336_(_1055_, _1052_, addr_tag[0]);
    or _1337_(_0191_, _1055_, _1054_);
    and _1338_(_1056_, _1053_, \cache_tags[6][1]);
    and _1339_(_1057_, _1052_, addr_tag[1]);
    or _1340_(_0192_, _1057_, _1056_);
    and _1341_(_1058_, _1053_, \cache_tags[6][2]);
    and _1342_(_1059_, _1052_, addr_tag[2]);
    or _1343_(_0193_, _1059_, _1058_);
    and _1344_(_1060_, _1053_, \cache_tags[6][3]);
    and _1345_(_1061_, _1052_, addr_tag[3]);
    or _1346_(_0194_, _1061_, _1060_);
    nor _1347_(_1062_, _1045_, cache_state[0]);
    and _1348_(_1063_, _1062_, _1044_);
    nor _1349_(_1064_, cache_state[1], cache_state[0]);
    and _1350_(_1065_, _1064_, _1044_);
    nor _1351_(_1066_, _1065_, _1063_);
    and _1352_(_1067_, _1066_, cache_ready);
    and _1353_(_1068_, _1062_, _1044_);
    or _1354_(_0195_, _1068_, _1067_);
    not _1355_(_1069_, cache_state[0]);
    nor _1356_(_1070_, cache_read, cache_write);
    and _1357_(_1071_, _1070_, _1047_);
    and _1358_(_1072_, _1070_, _1065_);
    nor _1359_(_1073_, _1072_, _1071_);
    nor _1360_(_1074_, _1073_, _1069_);
    not _1361_(_1075_, _1070_);
    and _1362_(_1076_, _1075_, _1065_);
    or _1363_(_1077_, _1065_, _1047_);
    and _1364_(_1078_, _1077_, _1076_);
    and _1365_(_1079_, _1078_, _1073_);
    or _1366_(_0196_, _1079_, _1074_);
    nor _1367_(_1080_, _1073_, _1045_);
    or _1368_(_1081_, cache_read, cache_write);
    and _1369_(_1082_, _1081_, _1047_);
    and _1370_(_1083_, _1082_, _1077_);
    and _1371_(_1084_, _1083_, _1073_);
    or _1372_(_0197_, _1084_, _1080_);
    nor _1373_(_0198_, _1073_, _1044_);
    nor _1374_(_1085_, _1076_, _1049_);
    and _1375_(_1086_, _1076_, addr_index[0]);
    or _1376_(_0199_, _1086_, _1085_);
    not _1377_(_1087_, access_index[1]);
    nor _1378_(_1088_, _1076_, _1087_);
    and _1379_(_1089_, _1076_, addr_index[1]);
    or _1380_(_0200_, _1089_, _1088_);
    not _1381_(_1090_, access_index[2]);
    nor _1382_(_1091_, _1076_, _1090_);
    and _1383_(_1092_, _1076_, addr_index[2]);
    or _1384_(_0201_, _1092_, _1091_);
    and _1385_(_1093_, _1087_, access_index[0]);
    and _1386_(_1094_, _1093_, _1090_);
    and _1387_(_1095_, _1094_, _1048_);
    not _1388_(_1096_, _1095_);
    and _1389_(_1097_, _1096_, \cache_data[1][0]);
    and _1390_(_1098_, _1095_, write_data[0]);
    or _1391_(_0202_, _1098_, _1097_);
    and _1392_(_1099_, _1096_, \cache_data[1][1]);
    and _1393_(_1100_, _1095_, write_data[1]);
    or _1394_(_0203_, _1100_, _1099_);
    and _1395_(_1101_, _1096_, \cache_data[1][2]);
    and _1396_(_1102_, _1095_, write_data[2]);
    or _1397_(_0204_, _1102_, _1101_);
    and _1398_(_1103_, _1096_, \cache_data[1][3]);
    and _1399_(_1104_, _1095_, write_data[3]);
    or _1400_(_0205_, _1104_, _1103_);
    and _1401_(_1105_, _1096_, \cache_data[1][4]);
    and _1402_(_1106_, _1095_, write_data[4]);
    or _1403_(_0206_, _1106_, _1105_);
    and _1404_(_1107_, _1096_, \cache_data[1][5]);
    and _1405_(_1108_, _1095_, write_data[5]);
    or _1406_(_0207_, _1108_, _1107_);
    and _1407_(_1109_, _1096_, \cache_data[1][6]);
    and _1408_(_1110_, _1095_, write_data[6]);
    or _1409_(_0208_, _1110_, _1109_);
    and _1410_(_1111_, _1096_, \cache_data[1][7]);
    and _1411_(_1112_, _1095_, write_data[7]);
    or _1412_(_0209_, _1112_, _1111_);
    and _1413_(_1113_, _1096_, \cache_data[1][8]);
    and _1414_(_1114_, _1095_, write_data[8]);
    or _1415_(_0210_, _1114_, _1113_);
    and _1416_(_1115_, _1096_, \cache_data[1][9]);
    and _1417_(_1116_, _1095_, write_data[9]);
    or _1418_(_0211_, _1116_, _1115_);
    and _1419_(_1117_, _1096_, \cache_data[1][10]);
    and _1420_(_1118_, _1095_, write_data[10]);
    or _1421_(_0212_, _1118_, _1117_);
    and _1422_(_1119_, _1096_, \cache_data[1][11]);
    and _1423_(_1120_, _1095_, write_data[11]);
    or _1424_(_0213_, _1120_, _1119_);
    and _1425_(_1121_, _1096_, \cache_data[1][12]);
    and _1426_(_1122_, _1095_, write_data[12]);
    or _1427_(_0214_, _1122_, _1121_);
    and _1428_(_1123_, _1096_, \cache_data[1][13]);
    and _1429_(_1124_, _1095_, write_data[13]);
    or _1430_(_0215_, _1124_, _1123_);
    and _1431_(_1125_, _1096_, \cache_data[1][14]);
    and _1432_(_1126_, _1095_, write_data[14]);
    or _1433_(_0216_, _1126_, _1125_);
    and _1434_(_1127_, _1096_, \cache_data[1][15]);
    and _1435_(_1128_, _1095_, write_data[15]);
    or _1436_(_0217_, _1128_, _1127_);
    and _1437_(_1129_, _1050_, _1090_);
    and _1438_(_1130_, _1129_, _1048_);
    not _1439_(_1131_, _1130_);
    and _1440_(_1132_, _1131_, \cache_data[2][0]);
    and _1441_(_1133_, _1130_, write_data[0]);
    or _1442_(_0218_, _1133_, _1132_);
    and _1443_(_1134_, _1131_, \cache_data[2][1]);
    and _1444_(_1135_, _1130_, write_data[1]);
    or _1445_(_0219_, _1135_, _1134_);
    and _1446_(_1136_, _1131_, \cache_data[2][2]);
    and _1447_(_1137_, _1130_, write_data[2]);
    or _1448_(_0220_, _1137_, _1136_);
    and _1449_(_1138_, _1131_, \cache_data[2][3]);
    and _1450_(_1139_, _1130_, write_data[3]);
    or _1451_(_0221_, _1139_, _1138_);
    and _1452_(_1140_, _1131_, \cache_data[2][4]);
    and _1453_(_1141_, _1130_, write_data[4]);
    or _1454_(_0222_, _1141_, _1140_);
    and _1455_(_1142_, _1131_, \cache_data[2][5]);
    and _1456_(_1143_, _1130_, write_data[5]);
    or _1457_(_0223_, _1143_, _1142_);
    and _1458_(_1144_, _1131_, \cache_data[2][6]);
    and _1459_(_1145_, _1130_, write_data[6]);
    or _1460_(_0224_, _1145_, _1144_);
    and _1461_(_1146_, _1131_, \cache_data[2][7]);
    and _1462_(_1147_, _1130_, write_data[7]);
    or _1463_(_0225_, _1147_, _1146_);
    and _1464_(_1148_, _1131_, \cache_data[2][8]);
    and _1465_(_1149_, _1130_, write_data[8]);
    or _1466_(_0226_, _1149_, _1148_);
    and _1467_(_1150_, _1131_, \cache_data[2][9]);
    and _1468_(_1151_, _1130_, write_data[9]);
    or _1469_(_0227_, _1151_, _1150_);
    and _1470_(_1152_, _1131_, \cache_data[2][10]);
    and _1471_(_1153_, _1130_, write_data[10]);
    or _1472_(_0228_, _1153_, _1152_);
    and _1473_(_1154_, _1131_, \cache_data[2][11]);
    and _1474_(_1155_, _1130_, write_data[11]);
    or _1475_(_0229_, _1155_, _1154_);
    and _1476_(_1156_, _1131_, \cache_data[2][12]);
    and _1477_(_1157_, _1130_, write_data[12]);
    or _1478_(_0230_, _1157_, _1156_);
    and _1479_(_1158_, _1131_, \cache_data[2][13]);
    and _1480_(_1159_, _1130_, write_data[13]);
    or _1481_(_0231_, _1159_, _1158_);
    and _1482_(_1160_, _1131_, \cache_data[2][14]);
    and _1483_(_1161_, _1130_, write_data[14]);
    or _1484_(_0232_, _1161_, _1160_);
    and _1485_(_1162_, _1131_, \cache_data[2][15]);
    and _1486_(_1163_, _1130_, write_data[15]);
    or _1487_(_0233_, _1163_, _1162_);
    nor _1488_(_1164_, access_index[1], access_index[0]);
    and _1489_(_1165_, _1164_, access_index[2]);
    and _1490_(_1166_, _1165_, _1048_);
    not _1491_(_1167_, _1166_);
    and _1492_(_1168_, _1167_, \cache_data[4][0]);
    and _1493_(_1169_, _1166_, write_data[0]);
    or _1494_(_0234_, _1169_, _1168_);
    and _1495_(_1170_, _1167_, \cache_data[4][1]);
    and _1496_(_1171_, _1166_, write_data[1]);
    or _1497_(_0235_, _1171_, _1170_);
    and _1498_(_1172_, _1167_, \cache_data[4][2]);
    and _1499_(_1173_, _1166_, write_data[2]);
    or _1500_(_0236_, _1173_, _1172_);
    and _1501_(_1174_, _1167_, \cache_data[4][3]);
    and _1502_(_1175_, _1166_, write_data[3]);
    or _1503_(_0237_, _1175_, _1174_);
    and _1504_(_1176_, _1167_, \cache_data[4][4]);
    and _1505_(_1177_, _1166_, write_data[4]);
    or _1506_(_0238_, _1177_, _1176_);
    and _1507_(_1178_, _1167_, \cache_data[4][5]);
    and _1508_(_1179_, _1166_, write_data[5]);
    or _1509_(_0239_, _1179_, _1178_);
    and _1510_(_1180_, _1167_, \cache_data[4][6]);
    and _1511_(_1181_, _1166_, write_data[6]);
    or _1512_(_0240_, _1181_, _1180_);
    and _1513_(_1182_, _1167_, \cache_data[4][7]);
    and _1514_(_1183_, _1166_, write_data[7]);
    or _1515_(_0241_, _1183_, _1182_);
    and _1516_(_1184_, _1167_, \cache_data[4][8]);
    and _1517_(_1185_, _1166_, write_data[8]);
    or _1518_(_0242_, _1185_, _1184_);
    and _1519_(_1186_, _1167_, \cache_data[4][9]);
    and _1520_(_1187_, _1166_, write_data[9]);
    or _1521_(_0243_, _1187_, _1186_);
    and _1522_(_1188_, _1167_, \cache_data[4][10]);
    and _1523_(_1189_, _1166_, write_data[10]);
    or _1524_(_0244_, _1189_, _1188_);
    and _1525_(_1190_, _1167_, \cache_data[4][11]);
    and _1526_(_1191_, _1166_, write_data[11]);
    or _1527_(_0245_, _1191_, _1190_);
    and _1528_(_1192_, _1167_, \cache_data[4][12]);
    and _1529_(_1193_, _1166_, write_data[12]);
    or _1530_(_0246_, _1193_, _1192_);
    and _1531_(_1194_, _1167_, \cache_data[4][13]);
    and _1532_(_1195_, _1166_, write_data[13]);
    or _1533_(_0247_, _1195_, _1194_);
    and _1534_(_1196_, _1167_, \cache_data[4][14]);
    and _1535_(_1197_, _1166_, write_data[14]);
    or _1536_(_0248_, _1197_, _1196_);
    and _1537_(_1198_, _1167_, \cache_data[4][15]);
    and _1538_(_1199_, _1166_, write_data[15]);
    or _1539_(_0249_, _1199_, _1198_);
    and _1540_(_1200_, _1093_, access_index[2]);
    and _1541_(_1201_, _1200_, _1048_);
    not _1542_(_1202_, _1201_);
    and _1543_(_1203_, _1202_, \cache_data[5][0]);
    and _1544_(_1204_, _1201_, write_data[0]);
    or _1545_(_0250_, _1204_, _1203_);
    and _1546_(_1205_, _1202_, \cache_data[5][1]);
    and _1547_(_1206_, _1201_, write_data[1]);
    or _1548_(_0251_, _1206_, _1205_);
    and _1549_(_1207_, _1202_, \cache_data[5][2]);
    and _1550_(_1208_, _1201_, write_data[2]);
    or _1551_(_0252_, _1208_, _1207_);
    and _1552_(_1209_, _1202_, \cache_data[5][3]);
    and _1553_(_1210_, _1201_, write_data[3]);
    or _1554_(_0253_, _1210_, _1209_);
    and _1555_(_1211_, _1202_, \cache_data[5][4]);
    and _1556_(_1212_, _1201_, write_data[4]);
    or _1557_(_0254_, _1212_, _1211_);
    and _1558_(_1213_, _1202_, \cache_data[5][5]);
    and _1559_(_1214_, _1201_, write_data[5]);
    or _1560_(_0255_, _1214_, _1213_);
    and _1561_(_1215_, _1202_, \cache_data[5][6]);
    and _1562_(_1216_, _1201_, write_data[6]);
    or _1563_(_0256_, _1216_, _1215_);
    and _1564_(_1217_, _1202_, \cache_data[5][7]);
    and _1565_(_1218_, _1201_, write_data[7]);
    or _1566_(_0257_, _1218_, _1217_);
    and _1567_(_1219_, _1202_, \cache_data[5][8]);
    and _1568_(_1220_, _1201_, write_data[8]);
    or _1569_(_0258_, _1220_, _1219_);
    and _1570_(_1221_, _1202_, \cache_data[5][9]);
    and _1571_(_1222_, _1201_, write_data[9]);
    or _1572_(_0259_, _1222_, _1221_);
    and _1573_(_1223_, _1202_, \cache_data[5][10]);
    and _1574_(_1224_, _1201_, write_data[10]);
    or _1575_(_0260_, _1224_, _1223_);
    and _1576_(_1225_, _1202_, \cache_data[5][11]);
    and _1577_(_1226_, _1201_, write_data[11]);
    or _1578_(_0261_, _1226_, _1225_);
    and _1579_(_1227_, _1202_, \cache_data[5][12]);
    and _1580_(_1228_, _1201_, write_data[12]);
    or _1581_(_0262_, _1228_, _1227_);
    and _1582_(_1229_, _1202_, \cache_data[5][13]);
    and _1583_(_1230_, _1201_, write_data[13]);
    or _1584_(_0263_, _1230_, _1229_);
    and _1585_(_1231_, _1202_, \cache_data[5][14]);
    and _1586_(_1232_, _1201_, write_data[14]);
    or _1587_(_0264_, _1232_, _1231_);
    and _1588_(_1233_, _1202_, \cache_data[5][15]);
    and _1589_(_1234_, _1201_, write_data[15]);
    or _1590_(_0265_, _1234_, _1233_);
    and _1591_(_1235_, _1053_, \cache_data[6][0]);
    and _1592_(_1236_, _1052_, write_data[0]);
    or _1593_(_0266_, _1236_, _1235_);
    and _1594_(_1237_, _1053_, \cache_data[6][1]);
    and _1595_(_1238_, _1052_, write_data[1]);
    or _1596_(_0267_, _1238_, _1237_);
    and _1597_(_1239_, _1053_, \cache_data[6][2]);
    and _1598_(_1240_, _1052_, write_data[2]);
    or _1599_(_0268_, _1240_, _1239_);
    and _1600_(_1241_, _1053_, \cache_data[6][3]);
    and _1601_(_1242_, _1052_, write_data[3]);
    or _1602_(_0269_, _1242_, _1241_);
    and _1603_(_1243_, _1053_, \cache_data[6][4]);
    and _1604_(_1244_, _1052_, write_data[4]);
    or _1605_(_0270_, _1244_, _1243_);
    and _1606_(_1245_, _1053_, \cache_data[6][5]);
    and _1607_(_1246_, _1052_, write_data[5]);
    or _1608_(_0271_, _1246_, _1245_);
    and _1609_(_1247_, _1053_, \cache_data[6][6]);
    and _1610_(_1248_, _1052_, write_data[6]);
    or _1611_(_0272_, _1248_, _1247_);
    and _1612_(_1249_, _1053_, \cache_data[6][7]);
    and _1613_(_1250_, _1052_, write_data[7]);
    or _1614_(_0273_, _1250_, _1249_);
    and _1615_(_1251_, _1053_, \cache_data[6][8]);
    and _1616_(_1252_, _1052_, write_data[8]);
    or _1617_(_0274_, _1252_, _1251_);
    and _1618_(_1253_, _1053_, \cache_data[6][9]);
    and _1619_(_1254_, _1052_, write_data[9]);
    or _1620_(_0275_, _1254_, _1253_);
    and _1621_(_1255_, _1053_, \cache_data[6][10]);
    and _1622_(_1256_, _1052_, write_data[10]);
    or _1623_(_0276_, _1256_, _1255_);
    and _1624_(_1257_, _1053_, \cache_data[6][11]);
    and _1625_(_1258_, _1052_, write_data[11]);
    or _1626_(_0277_, _1258_, _1257_);
    and _1627_(_1259_, _1053_, \cache_data[6][12]);
    and _1628_(_1260_, _1052_, write_data[12]);
    or _1629_(_0278_, _1260_, _1259_);
    and _1630_(_1261_, _1053_, \cache_data[6][13]);
    and _1631_(_1262_, _1052_, write_data[13]);
    or _1632_(_0279_, _1262_, _1261_);
    and _1633_(_1263_, _1053_, \cache_data[6][14]);
    and _1634_(_1264_, _1052_, write_data[14]);
    or _1635_(_0280_, _1264_, _1263_);
    and _1636_(_1265_, _1053_, \cache_data[6][15]);
    and _1637_(_1266_, _1052_, write_data[15]);
    or _1638_(_0281_, _1266_, _1265_);
    and _1639_(_1267_, access_index[1], access_index[0]);
    and _1640_(_1268_, _1267_, access_index[2]);
    and _1641_(_1269_, _1268_, _1048_);
    not _1642_(_1270_, _1269_);
    and _1643_(_1271_, _1270_, \cache_data[7][0]);
    and _1644_(_1272_, _1269_, write_data[0]);
    or _1645_(_0282_, _1272_, _1271_);
    and _1646_(_1273_, _1270_, \cache_data[7][1]);
    and _1647_(_1274_, _1269_, write_data[1]);
    or _1648_(_0283_, _1274_, _1273_);
    and _1649_(_1275_, _1270_, \cache_data[7][2]);
    and _1650_(_1276_, _1269_, write_data[2]);
    or _1651_(_0284_, _1276_, _1275_);
    and _1652_(_1277_, _1270_, \cache_data[7][3]);
    and _1653_(_1278_, _1269_, write_data[3]);
    or _1654_(_0285_, _1278_, _1277_);
    and _1655_(_1279_, _1270_, \cache_data[7][4]);
    and _1656_(_1280_, _1269_, write_data[4]);
    or _1657_(_0286_, _1280_, _1279_);
    and _1658_(_1281_, _1270_, \cache_data[7][5]);
    and _1659_(_1282_, _1269_, write_data[5]);
    or _1660_(_0287_, _1282_, _1281_);
    and _1661_(_1283_, _1270_, \cache_data[7][6]);
    and _1662_(_1284_, _1269_, write_data[6]);
    or _1663_(_0288_, _1284_, _1283_);
    and _1664_(_1285_, _1270_, \cache_data[7][7]);
    and _1665_(_1286_, _1269_, write_data[7]);
    or _1666_(_0289_, _1286_, _1285_);
    and _1667_(_1287_, _1270_, \cache_data[7][8]);
    and _1668_(_1288_, _1269_, write_data[8]);
    or _1669_(_0290_, _1288_, _1287_);
    and _1670_(_1289_, _1270_, \cache_data[7][9]);
    and _1671_(_1290_, _1269_, write_data[9]);
    or _1672_(_0291_, _1290_, _1289_);
    and _1673_(_1291_, _1270_, \cache_data[7][10]);
    and _1674_(_1292_, _1269_, write_data[10]);
    or _1675_(_0292_, _1292_, _1291_);
    and _1676_(_1293_, _1270_, \cache_data[7][11]);
    and _1677_(_1294_, _1269_, write_data[11]);
    or _1678_(_0293_, _1294_, _1293_);
    and _1679_(_1295_, _1270_, \cache_data[7][12]);
    and _1680_(_1296_, _1269_, write_data[12]);
    or _1681_(_0294_, _1296_, _1295_);
    and _1682_(_1297_, _1270_, \cache_data[7][13]);
    and _1683_(_1298_, _1269_, write_data[13]);
    or _1684_(_0295_, _1298_, _1297_);
    and _1685_(_1299_, _1270_, \cache_data[7][14]);
    and _1686_(_1300_, _1269_, write_data[14]);
    or _1687_(_0296_, _1300_, _1299_);
    and _1688_(_1301_, _1270_, \cache_data[7][15]);
    and _1689_(_1302_, _1269_, write_data[15]);
    or _1690_(_0297_, _1302_, _1301_);
    and _1691_(_1303_, _1164_, _1090_);
    and _1692_(_1304_, _1303_, _1048_);
    not _1693_(_1305_, _1304_);
    and _1694_(_1306_, _1305_, \cache_tags[0][0]);
    and _1695_(_1307_, _1304_, addr_tag[0]);
    or _1696_(_0298_, _1307_, _1306_);
    and _1697_(_1308_, _1305_, \cache_tags[0][1]);
    and _1698_(_1309_, _1304_, addr_tag[1]);
    or _1699_(_0299_, _1309_, _1308_);
    and _1700_(_1310_, _1305_, \cache_tags[0][2]);
    and _1701_(_1311_, _1304_, addr_tag[2]);
    or _1702_(_0300_, _1311_, _1310_);
    and _1703_(_1312_, _1305_, \cache_tags[0][3]);
    and _1704_(_1313_, _1304_, addr_tag[3]);
    or _1705_(_0301_, _1313_, _1312_);
    and _1706_(_1314_, _1096_, \cache_tags[1][0]);
    and _1707_(_1315_, _1095_, addr_tag[0]);
    or _1708_(_0302_, _1315_, _1314_);
    and _1709_(_1316_, _1096_, \cache_tags[1][1]);
    and _1710_(_1317_, _1095_, addr_tag[1]);
    or _1711_(_0303_, _1317_, _1316_);
    and _1712_(_1318_, _1096_, \cache_tags[1][2]);
    and _1713_(_1319_, _1095_, addr_tag[2]);
    or _1714_(_0304_, _1319_, _1318_);
    and _1715_(_1320_, _1096_, \cache_tags[1][3]);
    and _1716_(_1321_, _1095_, addr_tag[3]);
    or _1717_(_0305_, _1321_, _1320_);
    and _1718_(_1322_, _1131_, \cache_tags[2][0]);
    and _1719_(_1323_, _1130_, addr_tag[0]);
    or _1720_(_0306_, _1323_, _1322_);
    and _1721_(_0382_, _1131_, \cache_tags[2][1]);
    and _1722_(_0383_, _1130_, addr_tag[1]);
    or _1723_(_0307_, _0383_, _0382_);
    and _1724_(_0384_, _1131_, \cache_tags[2][2]);
    and _1725_(_0385_, _1130_, addr_tag[2]);
    or _1726_(_0308_, _0385_, _0384_);
    and _1727_(_0386_, _1131_, \cache_tags[2][3]);
    and _1728_(_0387_, _1130_, addr_tag[3]);
    or _1729_(_0309_, _0387_, _0386_);
    and _1730_(_0388_, _1267_, _1090_);
    and _1731_(_0389_, _0388_, _1048_);
    not _1732_(_0390_, _0389_);
    and _1733_(_0391_, _0390_, \cache_tags[3][0]);
    and _1734_(_0392_, _0389_, addr_tag[0]);
    or _1735_(_0310_, _0392_, _0391_);
    and _1736_(_0393_, _0390_, \cache_tags[3][1]);
    and _1737_(_0394_, _0389_, addr_tag[1]);
    or _1738_(_0311_, _0394_, _0393_);
    and _1739_(_0395_, _0390_, \cache_tags[3][2]);
    and _1740_(_0396_, _0389_, addr_tag[2]);
    or _1741_(_0312_, _0396_, _0395_);
    and _1742_(_0397_, _0390_, \cache_tags[3][3]);
    and _1743_(_0398_, _0389_, addr_tag[3]);
    or _1744_(_0313_, _0398_, _0397_);
    and _1745_(_0399_, _1167_, \cache_tags[4][0]);
    and _1746_(_0400_, _1166_, addr_tag[0]);
    or _1747_(_0314_, _0400_, _0399_);
    and _1748_(_0401_, _1167_, \cache_tags[4][1]);
    and _1749_(_0402_, _1166_, addr_tag[1]);
    or _1750_(_0315_, _0402_, _0401_);
    and _1751_(_0403_, _1167_, \cache_tags[4][2]);
    and _1752_(_0404_, _1166_, addr_tag[2]);
    or _1753_(_0316_, _0404_, _0403_);
    and _1754_(_0405_, _1167_, \cache_tags[4][3]);
    and _1755_(_0406_, _1166_, addr_tag[3]);
    or _1756_(_0317_, _0406_, _0405_);
    and _1757_(_0407_, _1202_, \cache_tags[5][0]);
    and _1758_(_0408_, _1201_, addr_tag[0]);
    or _1759_(_0318_, _0408_, _0407_);
    and _1760_(_0409_, _1202_, \cache_tags[5][1]);
    and _1761_(_0410_, _1201_, addr_tag[1]);
    or _1762_(_0319_, _0410_, _0409_);
    and _1763_(_0411_, _1202_, \cache_tags[5][2]);
    and _1764_(_0412_, _1201_, addr_tag[2]);
    or _1765_(_0320_, _0412_, _0411_);
    and _1766_(_0413_, _1202_, \cache_tags[5][3]);
    and _1767_(_0414_, _1201_, addr_tag[3]);
    or _1768_(_0321_, _0414_, _0413_);
    not _1769_(_0415_, cache_write);
    and _1770_(_0416_, _1047_, cache_read);
    and _1771_(_0417_, _0416_, _0415_);
    not _1772_(_0418_, _0417_);
    and _1773_(_0419_, _0418_, read_data[0]);
    nor _1774_(_0420_, addr_index[5], addr_index[4]);
    or _1775_(_0421_, addr_index[5], addr_index[4]);
    nand _1776_(_0422_, addr_index[3], addr_index[2]);
    not _1777_(_0423_, addr_index[2]);
    nand _1778_(_0424_, addr_index[3], _0423_);
    and _1779_(_0425_, _0424_, _0422_);
    or _1780_(_0426_, _0425_, _0421_);
    and _1781_(_0427_, _0426_, _0420_);
    not _1782_(_0428_, addr_index[1]);
    not _1783_(_0429_, addr_index[0]);
    and _1784_(_0430_, valid_bits[0], _0429_);
    and _1785_(_0431_, valid_bits[1], addr_index[0]);
    or _1786_(_0432_, _0431_, _0430_);
    and _1787_(_0433_, _0432_, _0428_);
    and _1788_(_0434_, valid_bits[2], _0429_);
    and _1789_(_0435_, valid_bits[3], addr_index[0]);
    or _1790_(_0436_, _0435_, _0434_);
    and _1791_(_0437_, _0436_, addr_index[1]);
    or _1792_(_0438_, _0437_, _0433_);
    and _1793_(_0439_, _0438_, _0423_);
    and _1794_(_0440_, valid_bits[4], _0429_);
    and _1795_(_0441_, valid_bits[5], addr_index[0]);
    or _1796_(_0442_, _0441_, _0440_);
    and _1797_(_0443_, _0442_, _0428_);
    and _1798_(_0444_, valid_bits[6], _0429_);
    and _1799_(_0445_, valid_bits[7], addr_index[0]);
    or _1800_(_0446_, _0445_, _0444_);
    and _1801_(_0447_, _0446_, addr_index[1]);
    or _1802_(_0448_, _0447_, _0443_);
    and _1803_(_0449_, _0448_, addr_index[2]);
    or _1804_(_0450_, _0449_, _0439_);
    and _1805_(_0451_, addr_index[1], addr_index[0]);
    and _1806_(_0452_, _0451_, addr_index[2]);
    and _1807_(_0453_, _0452_, \cache_tags[7][0]);
    and _1808_(_0454_, addr_index[1], _0429_);
    and _1809_(_0455_, _0454_, addr_index[2]);
    and _1810_(_0456_, _0455_, \cache_tags[6][0]);
    or _1811_(_0457_, _0456_, _0453_);
    and _1812_(_0458_, _0428_, addr_index[0]);
    and _1813_(_0459_, _0458_, addr_index[2]);
    and _1814_(_0460_, _0459_, \cache_tags[5][0]);
    nor _1815_(_0461_, addr_index[1], addr_index[0]);
    and _1816_(_0462_, _0461_, addr_index[2]);
    and _1817_(_0463_, _0462_, \cache_tags[4][0]);
    or _1818_(_0464_, _0463_, _0460_);
    or _1819_(_0465_, _0464_, _0457_);
    and _1820_(_0466_, _0451_, _0423_);
    and _1821_(_0467_, _0466_, \cache_tags[3][0]);
    and _1822_(_0468_, _0454_, _0423_);
    and _1823_(_0469_, _0468_, \cache_tags[2][0]);
    or _1824_(_0470_, _0469_, _0467_);
    and _1825_(_0471_, _0458_, _0423_);
    and _1826_(_0472_, _0471_, \cache_tags[1][0]);
    and _1827_(_0473_, _0461_, _0423_);
    and _1828_(_0474_, _0473_, \cache_tags[0][0]);
    or _1829_(_0475_, _0474_, _0472_);
    or _1830_(_0476_, _0475_, _0470_);
    or _1831_(_0477_, _0476_, _0465_);
    or _1832_(_0478_, _0455_, _0452_);
    or _1833_(_0479_, _0462_, _0459_);
    or _1834_(_0480_, _0479_, _0478_);
    or _1835_(_0481_, _0468_, _0466_);
    or _1836_(_0482_, _0473_, _0471_);
    or _1837_(_0483_, _0482_, _0481_);
    or _1838_(_0484_, _0483_, _0480_);
    and _1839_(_0485_, _0484_, _0477_);
    nand _1840_(_0486_, _0485_, _0427_);
    xor _1841_(_0487_, _0486_, addr_tag[0]);
    and _1842_(_0488_, _0452_, \cache_tags[7][1]);
    and _1843_(_0489_, _0455_, \cache_tags[6][1]);
    or _1844_(_0490_, _0489_, _0488_);
    and _1845_(_0491_, _0459_, \cache_tags[5][1]);
    and _1846_(_0492_, _0462_, \cache_tags[4][1]);
    or _1847_(_0493_, _0492_, _0491_);
    or _1848_(_0494_, _0493_, _0490_);
    and _1849_(_0495_, _0466_, \cache_tags[3][1]);
    and _1850_(_0496_, _0468_, \cache_tags[2][1]);
    or _1851_(_0497_, _0496_, _0495_);
    and _1852_(_0498_, _0471_, \cache_tags[1][1]);
    and _1853_(_0499_, _0473_, \cache_tags[0][1]);
    or _1854_(_0500_, _0499_, _0498_);
    or _1855_(_0501_, _0500_, _0497_);
    or _1856_(_0502_, _0501_, _0494_);
    and _1857_(_0503_, _0502_, _0484_);
    nand _1858_(_0504_, _0503_, _0427_);
    xor _1859_(_0505_, _0504_, addr_tag[1]);
    and _1860_(_0506_, _0505_, _0487_);
    and _1861_(_0507_, _0452_, \cache_tags[7][2]);
    and _1862_(_0508_, _0455_, \cache_tags[6][2]);
    or _1863_(_0509_, _0508_, _0507_);
    and _1864_(_0510_, _0459_, \cache_tags[5][2]);
    and _1865_(_0511_, _0462_, \cache_tags[4][2]);
    or _1866_(_0512_, _0511_, _0510_);
    or _1867_(_0513_, _0512_, _0509_);
    and _1868_(_0514_, _0466_, \cache_tags[3][2]);
    and _1869_(_0515_, _0468_, \cache_tags[2][2]);
    or _1870_(_0516_, _0515_, _0514_);
    and _1871_(_0517_, _0471_, \cache_tags[1][2]);
    and _1872_(_0518_, _0473_, \cache_tags[0][2]);
    or _1873_(_0519_, _0518_, _0517_);
    or _1874_(_0520_, _0519_, _0516_);
    or _1875_(_0521_, _0520_, _0513_);
    and _1876_(_0522_, _0521_, _0484_);
    nand _1877_(_0523_, _0522_, _0427_);
    xor _1878_(_0524_, _0523_, addr_tag[2]);
    and _1879_(_0525_, _0452_, \cache_tags[7][3]);
    and _1880_(_0526_, _0455_, \cache_tags[6][3]);
    or _1881_(_0527_, _0526_, _0525_);
    and _1882_(_0528_, _0459_, \cache_tags[5][3]);
    and _1883_(_0529_, _0462_, \cache_tags[4][3]);
    or _1884_(_0530_, _0529_, _0528_);
    or _1885_(_0531_, _0530_, _0527_);
    and _1886_(_0532_, _0466_, \cache_tags[3][3]);
    and _1887_(_0533_, _0468_, \cache_tags[2][3]);
    or _1888_(_0534_, _0533_, _0532_);
    and _1889_(_0535_, _0471_, \cache_tags[1][3]);
    and _1890_(_0536_, _0473_, \cache_tags[0][3]);
    or _1891_(_0537_, _0536_, _0535_);
    or _1892_(_0538_, _0537_, _0534_);
    or _1893_(_0539_, _0538_, _0531_);
    and _1894_(_0540_, _0539_, _0484_);
    nand _1895_(_0541_, _0540_, _0427_);
    xor _1896_(_0542_, _0541_, addr_tag[3]);
    and _1897_(_0543_, _0542_, _0524_);
    and _1898_(_0544_, _0543_, _0506_);
    and _1899_(_0545_, _0544_, _0450_);
    and _1900_(cache_hit, _0545_, _0427_);
    and _1901_(_0546_, _1268_, \cache_data[7][0]);
    and _1902_(_0547_, _1051_, \cache_data[6][0]);
    or _1903_(_0548_, _0547_, _0546_);
    and _1904_(_0549_, _1200_, \cache_data[5][0]);
    and _1905_(_0550_, _1165_, \cache_data[4][0]);
    or _1906_(_0551_, _0550_, _0549_);
    or _1907_(_0552_, _0551_, _0548_);
    and _1908_(_0553_, _0388_, \cache_data[3][0]);
    and _1909_(_0554_, _1129_, \cache_data[2][0]);
    or _1910_(_0555_, _0554_, _0553_);
    and _1911_(_0556_, _1094_, \cache_data[1][0]);
    and _1912_(_0557_, _1303_, \cache_data[0][0]);
    or _1913_(_0558_, _0557_, _0556_);
    or _1914_(_0559_, _0558_, _0555_);
    or _1915_(_0560_, _0559_, _0552_);
    or _1916_(_0561_, _1268_, _1051_);
    or _1917_(_0562_, _1200_, _1165_);
    or _1918_(_0563_, _0562_, _0561_);
    or _1919_(_0564_, _0388_, _1129_);
    or _1920_(_0565_, _1303_, _1094_);
    or _1921_(_0566_, _0565_, _0564_);
    or _1922_(_0567_, _0566_, _0563_);
    and _1923_(_0568_, _0567_, _0560_);
    and _1924_(_0569_, _0568_, cache_hit);
    and _1925_(_0570_, _0569_, cache_read);
    and _1926_(_0571_, _0570_, _0415_);
    and _1927_(_0572_, _0571_, _1047_);
    and _1928_(_0573_, _0572_, cache_hit);
    and _1929_(_0574_, _0573_, _0417_);
    or _1930_(_0322_, _0574_, _0419_);
    and _1931_(_0575_, _0418_, read_data[1]);
    and _1932_(_0576_, _1268_, \cache_data[7][1]);
    and _1933_(_0577_, _1051_, \cache_data[6][1]);
    or _1934_(_0578_, _0577_, _0576_);
    and _1935_(_0579_, _1200_, \cache_data[5][1]);
    and _1936_(_0580_, _1165_, \cache_data[4][1]);
    or _1937_(_0581_, _0580_, _0579_);
    or _1938_(_0582_, _0581_, _0578_);
    and _1939_(_0583_, _0388_, \cache_data[3][1]);
    and _1940_(_0584_, _1129_, \cache_data[2][1]);
    or _1941_(_0585_, _0584_, _0583_);
    and _1942_(_0586_, _1094_, \cache_data[1][1]);
    and _1943_(_0587_, _1303_, \cache_data[0][1]);
    or _1944_(_0588_, _0587_, _0586_);
    or _1945_(_0589_, _0588_, _0585_);
    or _1946_(_0590_, _0589_, _0582_);
    and _1947_(_0591_, _0590_, _0567_);
    and _1948_(_0592_, _0591_, cache_hit);
    and _1949_(_0593_, _0592_, cache_read);
    and _1950_(_0594_, _0593_, _0415_);
    and _1951_(_0595_, _0594_, _1047_);
    and _1952_(_0596_, _0595_, cache_hit);
    and _1953_(_0597_, _0596_, _0417_);
    or _1954_(_0323_, _0597_, _0575_);
    and _1955_(_0598_, _0418_, read_data[2]);
    and _1956_(_0599_, _1268_, \cache_data[7][2]);
    and _1957_(_0600_, _1051_, \cache_data[6][2]);
    or _1958_(_0601_, _0600_, _0599_);
    and _1959_(_0602_, _1200_, \cache_data[5][2]);
    and _1960_(_0603_, _1165_, \cache_data[4][2]);
    or _1961_(_0604_, _0603_, _0602_);
    or _1962_(_0605_, _0604_, _0601_);
    and _1963_(_0606_, _0388_, \cache_data[3][2]);
    and _1964_(_0607_, _1129_, \cache_data[2][2]);
    or _1965_(_0608_, _0607_, _0606_);
    and _1966_(_0609_, _1094_, \cache_data[1][2]);
    and _1967_(_0610_, _1303_, \cache_data[0][2]);
    or _1968_(_0611_, _0610_, _0609_);
    or _1969_(_0612_, _0611_, _0608_);
    or _1970_(_0613_, _0612_, _0605_);
    and _1971_(_0614_, _0613_, _0567_);
    and _1972_(_0615_, _0614_, cache_hit);
    and _1973_(_0616_, _0615_, cache_read);
    and _1974_(_0617_, _0616_, _0415_);
    and _1975_(_0618_, _0617_, _1047_);
    and _1976_(_0619_, _0618_, cache_hit);
    and _1977_(_0620_, _0619_, _0417_);
    or _1978_(_0324_, _0620_, _0598_);
    and _1979_(_0621_, _0418_, read_data[3]);
    and _1980_(_0622_, _1268_, \cache_data[7][3]);
    and _1981_(_0623_, _1051_, \cache_data[6][3]);
    or _1982_(_0624_, _0623_, _0622_);
    and _1983_(_0625_, _1200_, \cache_data[5][3]);
    and _1984_(_0626_, _1165_, \cache_data[4][3]);
    or _1985_(_0627_, _0626_, _0625_);
    or _1986_(_0628_, _0627_, _0624_);
    and _1987_(_0629_, _0388_, \cache_data[3][3]);
    and _1988_(_0630_, _1129_, \cache_data[2][3]);
    or _1989_(_0631_, _0630_, _0629_);
    and _1990_(_0632_, _1094_, \cache_data[1][3]);
    and _1991_(_0633_, _1303_, \cache_data[0][3]);
    or _1992_(_0634_, _0633_, _0632_);
    or _1993_(_0635_, _0634_, _0631_);
    or _1994_(_0636_, _0635_, _0628_);
    and _1995_(_0637_, _0636_, _0567_);
    and _1996_(_0638_, _0637_, cache_hit);
    and _1997_(_0639_, _0638_, cache_read);
    and _1998_(_0640_, _0639_, _0415_);
    and _1999_(_0641_, _0640_, _1047_);
    and _2000_(_0642_, _0641_, cache_hit);
    and _2001_(_0643_, _0642_, _0417_);
    or _2002_(_0325_, _0643_, _0621_);
    and _2003_(_0644_, _0418_, read_data[4]);
    and _2004_(_0645_, _1268_, \cache_data[7][4]);
    and _2005_(_0646_, _1051_, \cache_data[6][4]);
    or _2006_(_0647_, _0646_, _0645_);
    and _2007_(_0648_, _1200_, \cache_data[5][4]);
    and _2008_(_0649_, _1165_, \cache_data[4][4]);
    or _2009_(_0650_, _0649_, _0648_);
    or _2010_(_0651_, _0650_, _0647_);
    and _2011_(_0652_, _0388_, \cache_data[3][4]);
    and _2012_(_0653_, _1129_, \cache_data[2][4]);
    or _2013_(_0654_, _0653_, _0652_);
    and _2014_(_0655_, _1094_, \cache_data[1][4]);
    and _2015_(_0656_, _1303_, \cache_data[0][4]);
    or _2016_(_0657_, _0656_, _0655_);
    or _2017_(_0658_, _0657_, _0654_);
    or _2018_(_0659_, _0658_, _0651_);
    and _2019_(_0660_, _0659_, _0567_);
    and _2020_(_0661_, _0660_, cache_hit);
    and _2021_(_0662_, _0661_, cache_read);
    and _2022_(_0663_, _0662_, _0415_);
    and _2023_(_0664_, _0663_, _1047_);
    and _2024_(_0665_, _0664_, cache_hit);
    and _2025_(_0666_, _0665_, _0417_);
    or _2026_(_0326_, _0666_, _0644_);
    and _2027_(_0667_, _0418_, read_data[5]);
    and _2028_(_0668_, _1268_, \cache_data[7][5]);
    and _2029_(_0669_, _1051_, \cache_data[6][5]);
    or _2030_(_0670_, _0669_, _0668_);
    and _2031_(_0671_, _1200_, \cache_data[5][5]);
    and _2032_(_0672_, _1165_, \cache_data[4][5]);
    or _2033_(_0673_, _0672_, _0671_);
    or _2034_(_0674_, _0673_, _0670_);
    and _2035_(_0675_, _0388_, \cache_data[3][5]);
    and _2036_(_0676_, _1129_, \cache_data[2][5]);
    or _2037_(_0677_, _0676_, _0675_);
    and _2038_(_0678_, _1094_, \cache_data[1][5]);
    and _2039_(_0679_, _1303_, \cache_data[0][5]);
    or _2040_(_0680_, _0679_, _0678_);
    or _2041_(_0681_, _0680_, _0677_);
    or _2042_(_0682_, _0681_, _0674_);
    and _2043_(_0683_, _0682_, _0567_);
    and _2044_(_0684_, _0683_, cache_hit);
    and _2045_(_0685_, _0684_, cache_read);
    and _2046_(_0686_, _0685_, _0415_);
    and _2047_(_0687_, _0686_, _1047_);
    and _2048_(_0688_, _0687_, cache_hit);
    and _2049_(_0689_, _0688_, _0417_);
    or _2050_(_0327_, _0689_, _0667_);
    and _2051_(_0690_, _0418_, read_data[6]);
    and _2052_(_0691_, _1268_, \cache_data[7][6]);
    and _2053_(_0692_, _1051_, \cache_data[6][6]);
    or _2054_(_0693_, _0692_, _0691_);
    and _2055_(_0694_, _1200_, \cache_data[5][6]);
    and _2056_(_0695_, _1165_, \cache_data[4][6]);
    or _2057_(_0696_, _0695_, _0694_);
    or _2058_(_0697_, _0696_, _0693_);
    and _2059_(_0698_, _0388_, \cache_data[3][6]);
    and _2060_(_0699_, _1129_, \cache_data[2][6]);
    or _2061_(_0700_, _0699_, _0698_);
    and _2062_(_0701_, _1094_, \cache_data[1][6]);
    and _2063_(_0702_, _1303_, \cache_data[0][6]);
    or _2064_(_0703_, _0702_, _0701_);
    or _2065_(_0704_, _0703_, _0700_);
    or _2066_(_0705_, _0704_, _0697_);
    and _2067_(_0706_, _0705_, _0567_);
    and _2068_(_0707_, _0706_, cache_hit);
    and _2069_(_0708_, _0707_, cache_read);
    and _2070_(_0709_, _0708_, _0415_);
    and _2071_(_0710_, _0709_, _1047_);
    and _2072_(_0711_, _0710_, cache_hit);
    and _2073_(_0712_, _0711_, _0417_);
    or _2074_(_0328_, _0712_, _0690_);
    and _2075_(_0713_, _0418_, read_data[7]);
    and _2076_(_0714_, _1268_, \cache_data[7][7]);
    and _2077_(_0715_, _1051_, \cache_data[6][7]);
    or _2078_(_0716_, _0715_, _0714_);
    and _2079_(_0717_, _1200_, \cache_data[5][7]);
    and _2080_(_0718_, _1165_, \cache_data[4][7]);
    or _2081_(_0719_, _0718_, _0717_);
    or _2082_(_0720_, _0719_, _0716_);
    and _2083_(_0721_, _0388_, \cache_data[3][7]);
    and _2084_(_0722_, _1129_, \cache_data[2][7]);
    or _2085_(_0723_, _0722_, _0721_);
    and _2086_(_0724_, _1094_, \cache_data[1][7]);
    and _2087_(_0725_, _1303_, \cache_data[0][7]);
    or _2088_(_0726_, _0725_, _0724_);
    or _2089_(_0727_, _0726_, _0723_);
    or _2090_(_0728_, _0727_, _0720_);
    and _2091_(_0729_, _0728_, _0567_);
    and _2092_(_0730_, _0729_, cache_hit);
    and _2093_(_0731_, _0730_, cache_read);
    and _2094_(_0732_, _0731_, _0415_);
    and _2095_(_0733_, _0732_, _1047_);
    and _2096_(_0734_, _0733_, cache_hit);
    and _2097_(_0735_, _0734_, _0417_);
    or _2098_(_0329_, _0735_, _0713_);
    and _2099_(_0736_, _0418_, read_data[8]);
    and _2100_(_0737_, _1268_, \cache_data[7][8]);
    and _2101_(_0738_, _1051_, \cache_data[6][8]);
    or _2102_(_0739_, _0738_, _0737_);
    and _2103_(_0740_, _1200_, \cache_data[5][8]);
    and _2104_(_0741_, _1165_, \cache_data[4][8]);
    or _2105_(_0742_, _0741_, _0740_);
    or _2106_(_0743_, _0742_, _0739_);
    and _2107_(_0744_, _0388_, \cache_data[3][8]);
    and _2108_(_0745_, _1129_, \cache_data[2][8]);
    or _2109_(_0746_, _0745_, _0744_);
    and _2110_(_0747_, _1094_, \cache_data[1][8]);
    and _2111_(_0748_, _1303_, \cache_data[0][8]);
    or _2112_(_0749_, _0748_, _0747_);
    or _2113_(_0750_, _0749_, _0746_);
    or _2114_(_0751_, _0750_, _0743_);
    and _2115_(_0752_, _0751_, _0567_);
    and _2116_(_0753_, _0752_, cache_hit);
    and _2117_(_0754_, _0753_, cache_read);
    and _2118_(_0755_, _0754_, _0415_);
    and _2119_(_0756_, _0755_, _1047_);
    and _2120_(_0757_, _0756_, cache_hit);
    and _2121_(_0758_, _0757_, _0417_);
    or _2122_(_0330_, _0758_, _0736_);
    and _2123_(_0759_, _0418_, read_data[9]);
    and _2124_(_0760_, _1268_, \cache_data[7][9]);
    and _2125_(_0761_, _1051_, \cache_data[6][9]);
    or _2126_(_0762_, _0761_, _0760_);
    and _2127_(_0763_, _1200_, \cache_data[5][9]);
    and _2128_(_0764_, _1165_, \cache_data[4][9]);
    or _2129_(_0765_, _0764_, _0763_);
    or _2130_(_0766_, _0765_, _0762_);
    and _2131_(_0767_, _0388_, \cache_data[3][9]);
    and _2132_(_0768_, _1129_, \cache_data[2][9]);
    or _2133_(_0769_, _0768_, _0767_);
    and _2134_(_0770_, _1094_, \cache_data[1][9]);
    and _2135_(_0771_, _1303_, \cache_data[0][9]);
    or _2136_(_0772_, _0771_, _0770_);
    or _2137_(_0773_, _0772_, _0769_);
    or _2138_(_0774_, _0773_, _0766_);
    and _2139_(_0775_, _0774_, _0567_);
    and _2140_(_0776_, _0775_, cache_hit);
    and _2141_(_0777_, _0776_, cache_read);
    and _2142_(_0778_, _0777_, _0415_);
    and _2143_(_0779_, _0778_, _1047_);
    and _2144_(_0780_, _0779_, cache_hit);
    and _2145_(_0781_, _0780_, _0417_);
    or _2146_(_0331_, _0781_, _0759_);
    and _2147_(_0782_, _0418_, read_data[10]);
    and _2148_(_0783_, _1268_, \cache_data[7][10]);
    and _2149_(_0784_, _1051_, \cache_data[6][10]);
    or _2150_(_0785_, _0784_, _0783_);
    and _2151_(_0786_, _1200_, \cache_data[5][10]);
    and _2152_(_0787_, _1165_, \cache_data[4][10]);
    or _2153_(_0788_, _0787_, _0786_);
    or _2154_(_0789_, _0788_, _0785_);
    and _2155_(_0790_, _0388_, \cache_data[3][10]);
    and _2156_(_0791_, _1129_, \cache_data[2][10]);
    or _2157_(_0792_, _0791_, _0790_);
    and _2158_(_0793_, _1094_, \cache_data[1][10]);
    and _2159_(_0794_, _1303_, \cache_data[0][10]);
    or _2160_(_0795_, _0794_, _0793_);
    or _2161_(_0796_, _0795_, _0792_);
    or _2162_(_0797_, _0796_, _0789_);
    and _2163_(_0798_, _0797_, _0567_);
    and _2164_(_0799_, _0798_, cache_hit);
    and _2165_(_0800_, _0799_, cache_read);
    and _2166_(_0801_, _0800_, _0415_);
    and _2167_(_0802_, _0801_, _1047_);
    and _2168_(_0803_, _0802_, cache_hit);
    and _2169_(_0804_, _0803_, _0417_);
    or _2170_(_0332_, _0804_, _0782_);
    and _2171_(_0805_, _0418_, read_data[11]);
    and _2172_(_0806_, _1268_, \cache_data[7][11]);
    and _2173_(_0807_, _1051_, \cache_data[6][11]);
    or _2174_(_0808_, _0807_, _0806_);
    and _2175_(_0809_, _1200_, \cache_data[5][11]);
    and _2176_(_0810_, _1165_, \cache_data[4][11]);
    or _2177_(_0811_, _0810_, _0809_);
    or _2178_(_0812_, _0811_, _0808_);
    and _2179_(_0813_, _0388_, \cache_data[3][11]);
    and _2180_(_0814_, _1129_, \cache_data[2][11]);
    or _2181_(_0815_, _0814_, _0813_);
    and _2182_(_0816_, _1094_, \cache_data[1][11]);
    and _2183_(_0817_, _1303_, \cache_data[0][11]);
    or _2184_(_0818_, _0817_, _0816_);
    or _2185_(_0819_, _0818_, _0815_);
    or _2186_(_0820_, _0819_, _0812_);
    and _2187_(_0821_, _0820_, _0567_);
    and _2188_(_0822_, _0821_, cache_hit);
    and _2189_(_0823_, _0822_, cache_read);
    and _2190_(_0824_, _0823_, _0415_);
    and _2191_(_0825_, _0824_, _1047_);
    and _2192_(_0826_, _0825_, cache_hit);
    and _2193_(_0827_, _0826_, _0417_);
    or _2194_(_0333_, _0827_, _0805_);
    and _2195_(_0828_, _0418_, read_data[12]);
    and _2196_(_0829_, _1268_, \cache_data[7][12]);
    and _2197_(_0830_, _1051_, \cache_data[6][12]);
    or _2198_(_0831_, _0830_, _0829_);
    and _2199_(_0832_, _1200_, \cache_data[5][12]);
    and _2200_(_0833_, _1165_, \cache_data[4][12]);
    or _2201_(_0834_, _0833_, _0832_);
    or _2202_(_0835_, _0834_, _0831_);
    and _2203_(_0836_, _0388_, \cache_data[3][12]);
    and _2204_(_0837_, _1129_, \cache_data[2][12]);
    or _2205_(_0838_, _0837_, _0836_);
    and _2206_(_0839_, _1094_, \cache_data[1][12]);
    and _2207_(_0840_, _1303_, \cache_data[0][12]);
    or _2208_(_0841_, _0840_, _0839_);
    or _2209_(_0842_, _0841_, _0838_);
    or _2210_(_0843_, _0842_, _0835_);
    and _2211_(_0844_, _0843_, _0567_);
    and _2212_(_0845_, _0844_, cache_hit);
    and _2213_(_0846_, _0845_, cache_read);
    and _2214_(_0847_, _0846_, _0415_);
    and _2215_(_0848_, _0847_, _1047_);
    and _2216_(_0849_, _0848_, cache_hit);
    and _2217_(_0850_, _0849_, _0417_);
    or _2218_(_0334_, _0850_, _0828_);
    and _2219_(_0851_, _0418_, read_data[13]);
    and _2220_(_0852_, _1268_, \cache_data[7][13]);
    and _2221_(_0853_, _1051_, \cache_data[6][13]);
    or _2222_(_0854_, _0853_, _0852_);
    and _2223_(_0855_, _1200_, \cache_data[5][13]);
    and _2224_(_0856_, _1165_, \cache_data[4][13]);
    or _2225_(_0857_, _0856_, _0855_);
    or _2226_(_0858_, _0857_, _0854_);
    and _2227_(_0859_, _0388_, \cache_data[3][13]);
    and _2228_(_0860_, _1129_, \cache_data[2][13]);
    or _2229_(_0861_, _0860_, _0859_);
    and _2230_(_0862_, _1094_, \cache_data[1][13]);
    and _2231_(_0863_, _1303_, \cache_data[0][13]);
    or _2232_(_0864_, _0863_, _0862_);
    or _2233_(_0865_, _0864_, _0861_);
    or _2234_(_0866_, _0865_, _0858_);
    and _2235_(_0867_, _0866_, _0567_);
    and _2236_(_0868_, _0867_, cache_hit);
    and _2237_(_0869_, _0868_, cache_read);
    and _2238_(_0870_, _0869_, _0415_);
    and _2239_(_0871_, _0870_, _1047_);
    and _2240_(_0872_, _0871_, cache_hit);
    and _2241_(_0873_, _0872_, _0417_);
    or _2242_(_0335_, _0873_, _0851_);
    and _2243_(_0874_, _0418_, read_data[14]);
    and _2244_(_0875_, _1268_, \cache_data[7][14]);
    and _2245_(_0876_, _1051_, \cache_data[6][14]);
    or _2246_(_0877_, _0876_, _0875_);
    and _2247_(_0878_, _1200_, \cache_data[5][14]);
    and _2248_(_0879_, _1165_, \cache_data[4][14]);
    or _2249_(_0880_, _0879_, _0878_);
    or _2250_(_0881_, _0880_, _0877_);
    and _2251_(_0882_, _0388_, \cache_data[3][14]);
    and _2252_(_0883_, _1129_, \cache_data[2][14]);
    or _2253_(_0884_, _0883_, _0882_);
    and _2254_(_0885_, _1094_, \cache_data[1][14]);
    and _2255_(_0886_, _1303_, \cache_data[0][14]);
    or _2256_(_0887_, _0886_, _0885_);
    or _2257_(_0888_, _0887_, _0884_);
    or _2258_(_0889_, _0888_, _0881_);
    and _2259_(_0890_, _0889_, _0567_);
    and _2260_(_0891_, _0890_, cache_hit);
    and _2261_(_0892_, _0891_, cache_read);
    and _2262_(_0893_, _0892_, _0415_);
    and _2263_(_0894_, _0893_, _1047_);
    and _2264_(_0895_, _0894_, cache_hit);
    and _2265_(_0896_, _0895_, _0417_);
    or _2266_(_0336_, _0896_, _0874_);
    and _2267_(_0897_, _0418_, read_data[15]);
    and _2268_(_0898_, _1268_, \cache_data[7][15]);
    and _2269_(_0899_, _1051_, \cache_data[6][15]);
    or _2270_(_0900_, _0899_, _0898_);
    and _2271_(_0901_, _1200_, \cache_data[5][15]);
    and _2272_(_0902_, _1165_, \cache_data[4][15]);
    or _2273_(_0903_, _0902_, _0901_);
    or _2274_(_0904_, _0903_, _0900_);
    and _2275_(_0905_, _0388_, \cache_data[3][15]);
    and _2276_(_0906_, _1129_, \cache_data[2][15]);
    or _2277_(_0907_, _0906_, _0905_);
    and _2278_(_0908_, _1094_, \cache_data[1][15]);
    and _2279_(_0909_, _1303_, \cache_data[0][15]);
    or _2280_(_0910_, _0909_, _0908_);
    or _2281_(_0911_, _0910_, _0907_);
    or _2282_(_0912_, _0911_, _0904_);
    and _2283_(_0913_, _0912_, _0567_);
    and _2284_(_0914_, _0913_, cache_hit);
    and _2285_(_0915_, _0914_, cache_read);
    and _2286_(_0916_, _0915_, _0415_);
    and _2287_(_0917_, _0916_, _1047_);
    and _2288_(_0918_, _0917_, cache_hit);
    and _2289_(_0919_, _0918_, _0417_);
    or _2290_(_0337_, _0919_, _0897_);
    and _2291_(_0920_, _1270_, \cache_tags[7][0]);
    and _2292_(_0921_, _1269_, addr_tag[0]);
    or _2293_(_0338_, _0921_, _0920_);
    and _2294_(_0922_, _1270_, \cache_tags[7][1]);
    and _2295_(_0923_, _1269_, addr_tag[1]);
    or _2296_(_0339_, _0923_, _0922_);
    and _2297_(_0924_, _1270_, \cache_tags[7][2]);
    and _2298_(_0925_, _1269_, addr_tag[2]);
    or _2299_(_0340_, _0925_, _0924_);
    and _2300_(_0926_, _1270_, \cache_tags[7][3]);
    and _2301_(_0927_, _1269_, addr_tag[3]);
    or _2302_(_0341_, _0927_, _0926_);
    and _2303_(_0928_, _0390_, \cache_data[3][0]);
    and _2304_(_0929_, _0389_, write_data[0]);
    or _2305_(_0342_, _0929_, _0928_);
    and _2306_(_0930_, _0390_, \cache_data[3][1]);
    and _2307_(_0931_, _0389_, write_data[1]);
    or _2308_(_0343_, _0931_, _0930_);
    and _2309_(_0932_, _0390_, \cache_data[3][2]);
    and _2310_(_0933_, _0389_, write_data[2]);
    or _2311_(_0344_, _0933_, _0932_);
    and _2312_(_0934_, _0390_, \cache_data[3][3]);
    and _2313_(_0935_, _0389_, write_data[3]);
    or _2314_(_0345_, _0935_, _0934_);
    and _2315_(_0936_, _0390_, \cache_data[3][4]);
    and _2316_(_0937_, _0389_, write_data[4]);
    or _2317_(_0346_, _0937_, _0936_);
    and _2318_(_0938_, _0390_, \cache_data[3][5]);
    and _2319_(_0939_, _0389_, write_data[5]);
    or _2320_(_0347_, _0939_, _0938_);
    and _2321_(_0940_, _0390_, \cache_data[3][6]);
    and _2322_(_0941_, _0389_, write_data[6]);
    or _2323_(_0348_, _0941_, _0940_);
    and _2324_(_0942_, _0390_, \cache_data[3][7]);
    and _2325_(_0943_, _0389_, write_data[7]);
    or _2326_(_0349_, _0943_, _0942_);
    and _2327_(_0944_, _0390_, \cache_data[3][8]);
    and _2328_(_0945_, _0389_, write_data[8]);
    or _2329_(_0350_, _0945_, _0944_);
    and _2330_(_0946_, _0390_, \cache_data[3][9]);
    and _2331_(_0947_, _0389_, write_data[9]);
    or _2332_(_0351_, _0947_, _0946_);
    and _2333_(_0948_, _0390_, \cache_data[3][10]);
    and _2334_(_0949_, _0389_, write_data[10]);
    or _2335_(_0352_, _0949_, _0948_);
    and _2336_(_0950_, _0390_, \cache_data[3][11]);
    and _2337_(_0951_, _0389_, write_data[11]);
    or _2338_(_0353_, _0951_, _0950_);
    and _2339_(_0952_, _0390_, \cache_data[3][12]);
    and _2340_(_0953_, _0389_, write_data[12]);
    or _2341_(_0354_, _0953_, _0952_);
    and _2342_(_0954_, _0390_, \cache_data[3][13]);
    and _2343_(_0955_, _0389_, write_data[13]);
    or _2344_(_0355_, _0955_, _0954_);
    and _2345_(_0956_, _0390_, \cache_data[3][14]);
    and _2346_(_0957_, _0389_, write_data[14]);
    or _2347_(_0356_, _0957_, _0956_);
    and _2348_(_0958_, _0390_, \cache_data[3][15]);
    and _2349_(_0959_, _0389_, write_data[15]);
    or _2350_(_0357_, _0959_, _0958_);
    and _2351_(_0960_, _1305_, \cache_data[0][0]);
    and _2352_(_0961_, _1304_, write_data[0]);
    or _2353_(_0358_, _0961_, _0960_);
    and _2354_(_0962_, _1305_, \cache_data[0][1]);
    and _2355_(_0963_, _1304_, write_data[1]);
    or _2356_(_0359_, _0963_, _0962_);
    and _2357_(_0964_, _1305_, \cache_data[0][2]);
    and _2358_(_0965_, _1304_, write_data[2]);
    or _2359_(_0360_, _0965_, _0964_);
    and _2360_(_0966_, _1305_, \cache_data[0][3]);
    and _2361_(_0967_, _1304_, write_data[3]);
    or _2362_(_0361_, _0967_, _0966_);
    and _2363_(_0968_, _1305_, \cache_data[0][4]);
    and _2364_(_0969_, _1304_, write_data[4]);
    or _2365_(_0362_, _0969_, _0968_);
    and _2366_(_0970_, _1305_, \cache_data[0][5]);
    and _2367_(_0971_, _1304_, write_data[5]);
    or _2368_(_0363_, _0971_, _0970_);
    and _2369_(_0972_, _1305_, \cache_data[0][6]);
    and _2370_(_0973_, _1304_, write_data[6]);
    or _2371_(_0364_, _0973_, _0972_);
    and _2372_(_0974_, _1305_, \cache_data[0][7]);
    and _2373_(_0975_, _1304_, write_data[7]);
    or _2374_(_0365_, _0975_, _0974_);
    and _2375_(_0976_, _1305_, \cache_data[0][8]);
    and _2376_(_0977_, _1304_, write_data[8]);
    or _2377_(_0366_, _0977_, _0976_);
    and _2378_(_0978_, _1305_, \cache_data[0][9]);
    and _2379_(_0979_, _1304_, write_data[9]);
    or _2380_(_0367_, _0979_, _0978_);
    and _2381_(_0980_, _1305_, \cache_data[0][10]);
    and _2382_(_0981_, _1304_, write_data[10]);
    or _2383_(_0368_, _0981_, _0980_);
    and _2384_(_0982_, _1305_, \cache_data[0][11]);
    and _2385_(_0983_, _1304_, write_data[11]);
    or _2386_(_0369_, _0983_, _0982_);
    and _2387_(_0984_, _1305_, \cache_data[0][12]);
    and _2388_(_0985_, _1304_, write_data[12]);
    or _2389_(_0370_, _0985_, _0984_);
    and _2390_(_0986_, _1305_, \cache_data[0][13]);
    and _2391_(_0987_, _1304_, write_data[13]);
    or _2392_(_0371_, _0987_, _0986_);
    and _2393_(_0988_, _1305_, \cache_data[0][14]);
    and _2394_(_0989_, _1304_, write_data[14]);
    or _2395_(_0372_, _0989_, _0988_);
    and _2396_(_0990_, _1305_, \cache_data[0][15]);
    and _2397_(_0991_, _1304_, write_data[15]);
    or _2398_(_0373_, _0991_, _0990_);
    not _2399_(_0992_, _1048_);
    and _2400_(_0993_, _0992_, valid_bits[0]);
    and _2401_(_0994_, _1303_, _1049_);
    xnor _2402_(_0995_, access_index[1], access_index[0]);
    and _2403_(_0996_, _0995_, _0994_);
    xor _2404_(_0997_, _1164_, access_index[2]);
    and _2405_(_0998_, _0997_, _0996_);
    and _2406_(_0999_, _0998_, _1303_);
    or _2407_(_1000_, _0999_, valid_bits[0]);
    and _2408_(_1001_, _1000_, _1048_);
    or _2409_(_0374_, _1001_, _0993_);
    and _2410_(_1002_, _0992_, valid_bits[1]);
    not _2411_(_1003_, _1303_);
    not _2412_(_1004_, _0997_);
    and _2413_(_1005_, _1087_, access_index[0]);
    and _2414_(_1006_, _1005_, _1004_);
    and _2415_(_1007_, _1006_, _1003_);
    or _2416_(_1008_, _1007_, valid_bits[1]);
    and _2417_(_1009_, _1008_, _1048_);
    or _2418_(_0375_, _1009_, _1002_);
    and _2419_(_1010_, _0992_, valid_bits[2]);
    and _2420_(_1011_, access_index[1], _1049_);
    and _2421_(_1012_, _1011_, _1004_);
    and _2422_(_1013_, _1012_, _1003_);
    or _2423_(_1014_, _1013_, valid_bits[2]);
    and _2424_(_1015_, _1014_, _1048_);
    or _2425_(_0376_, _1015_, _1010_);
    and _2426_(_1016_, _0992_, valid_bits[3]);
    and _2427_(_1017_, access_index[1], access_index[0]);
    and _2428_(_1018_, _1017_, _1004_);
    and _2429_(_1019_, _1018_, _1003_);
    or _2430_(_1020_, _1019_, valid_bits[3]);
    and _2431_(_1021_, _1020_, _1048_);
    or _2432_(_0377_, _1021_, _1016_);
    and _2433_(_1022_, _0992_, valid_bits[4]);
    nor _2434_(_1023_, _1303_, access_index[0]);
    and _2435_(_1024_, _1023_, _0995_);
    and _2436_(_1025_, _1024_, _1004_);
    and _2437_(_1026_, _1025_, _1003_);
    or _2438_(_1027_, _1026_, valid_bits[4]);
    and _2439_(_1028_, _1027_, _1048_);
    or _2440_(_0378_, _1028_, _1022_);
    and _2441_(_1029_, _0992_, valid_bits[5]);
    and _2442_(_1030_, _1005_, _0997_);
    and _2443_(_1031_, _1030_, _1003_);
    or _2444_(_1032_, _1031_, valid_bits[5]);
    and _2445_(_1033_, _1032_, _1048_);
    or _2446_(_0379_, _1033_, _1029_);
    and _2447_(_1034_, _0992_, valid_bits[6]);
    and _2448_(_1035_, _1011_, _0997_);
    and _2449_(_1036_, _1035_, _1003_);
    or _2450_(_1037_, _1036_, valid_bits[6]);
    and _2451_(_1038_, _1037_, _1048_);
    or _2452_(_0380_, _1038_, _1034_);
    and _2453_(_1039_, _0992_, valid_bits[7]);
    and _2454_(_1040_, _1017_, _0997_);
    and _2455_(_1041_, _1040_, _1003_);
    or _2456_(_1042_, _1041_, valid_bits[7]);
    and _2457_(_1043_, _1042_, _1048_);
    or _2458_(_0381_, _1043_, _1039_);
    not _2459_(_0001_, rst);
    not _2460_(_0002_, rst);
    not _2461_(_0003_, rst);
    not _2462_(_0004_, rst);
    not _2463_(_0005_, rst);
    not _2464_(_0006_, rst);
    not _2465_(_0007_, rst);
    not _2466_(_0008_, rst);
    not _2467_(_0009_, rst);
    not _2468_(_0010_, rst);
    not _2469_(_0011_, rst);
    not _2470_(_0012_, rst);
    not _2471_(_0013_, rst);
    not _2472_(_0014_, rst);
    not _2473_(_0015_, rst);
    not _2474_(_0016_, rst);
    not _2475_(_0017_, rst);
    not _2476_(_0018_, rst);
    not _2477_(_0019_, rst);
    not _2478_(_0020_, rst);
    not _2479_(_0021_, rst);
    not _2480_(_0022_, rst);
    not _2481_(_0023_, rst);
    not _2482_(_0024_, rst);
    not _2483_(_0025_, rst);
    not _2484_(_0026_, rst);
    not _2485_(_0027_, rst);
    not _2486_(_0028_, rst);
    not _2487_(_0029_, rst);
    not _2488_(_0030_, rst);
    not _2489_(_0031_, rst);
    not _2490_(_0032_, rst);
    not _2491_(_0033_, rst);
    not _2492_(_0034_, rst);
    not _2493_(_0035_, rst);
    not _2494_(_0036_, rst);
    not _2495_(_0037_, rst);
    not _2496_(_0038_, rst);
    not _2497_(_0039_, rst);
    not _2498_(_0040_, rst);
    not _2499_(_0041_, rst);
    not _2500_(_0042_, rst);
    not _2501_(_0043_, rst);
    not _2502_(_0044_, rst);
    not _2503_(_0045_, rst);
    not _2504_(_0046_, rst);
    not _2505_(_0047_, rst);
    not _2506_(_0048_, rst);
    not _2507_(_0049_, rst);
    not _2508_(_0050_, rst);
    not _2509_(_0051_, rst);
    not _2510_(_0052_, rst);
    not _2511_(_0053_, rst);
    not _2512_(_0054_, rst);
    not _2513_(_0055_, rst);
    not _2514_(_0056_, rst);
    not _2515_(_0057_, rst);
    not _2516_(_0058_, rst);
    not _2517_(_0059_, rst);
    not _2518_(_0060_, rst);
    not _2519_(_0061_, rst);
    not _2520_(_0062_, rst);
    not _2521_(_0063_, rst);
    not _2522_(_0064_, rst);
    not _2523_(_0065_, rst);
    not _2524_(_0066_, rst);
    not _2525_(_0067_, rst);
    not _2526_(_0068_, rst);
    not _2527_(_0069_, rst);
    not _2528_(_0070_, rst);
    not _2529_(_0071_, rst);
    not _2530_(_0072_, rst);
    not _2531_(_0073_, rst);
    not _2532_(_0074_, rst);
    not _2533_(_0075_, rst);
    not _2534_(_0076_, rst);
    not _2535_(_0077_, rst);
    not _2536_(_0078_, rst);
    not _2537_(_0079_, rst);
    not _2538_(_0080_, rst);
    not _2539_(_0081_, rst);
    not _2540_(_0082_, rst);
    not _2541_(_0083_, rst);
    not _2542_(_0084_, rst);
    not _2543_(_0085_, rst);
    not _2544_(_0086_, rst);
    not _2545_(_0087_, rst);
    not _2546_(_0088_, rst);
    not _2547_(_0089_, rst);
    not _2548_(_0090_, rst);
    not _2549_(_0091_, rst);
    not _2550_(_0092_, rst);
    not _2551_(_0093_, rst);
    not _2552_(_0094_, rst);
    not _2553_(_0095_, rst);
    not _2554_(_0096_, rst);
    not _2555_(_0097_, rst);
    not _2556_(_0098_, rst);
    not _2557_(_0099_, rst);
    not _2558_(_0100_, rst);
    not _2559_(_0101_, rst);
    not _2560_(_0102_, rst);
    not _2561_(_0103_, rst);
    not _2562_(_0104_, rst);
    not _2563_(_0105_, rst);
    not _2564_(_0106_, rst);
    not _2565_(_0107_, rst);
    not _2566_(_0108_, rst);
    not _2567_(_0109_, rst);
    not _2568_(_0110_, rst);
    not _2569_(_0111_, rst);
    not _2570_(_0112_, rst);
    not _2571_(_0113_, rst);
    not _2572_(_0114_, rst);
    not _2573_(_0115_, rst);
    not _2574_(_0116_, rst);
    not _2575_(_0117_, rst);
    not _2576_(_0118_, rst);
    not _2577_(_0119_, rst);
    not _2578_(_0120_, rst);
    not _2579_(_0121_, rst);
    not _2580_(_0122_, rst);
    not _2581_(_0123_, rst);
    not _2582_(_0124_, rst);
    not _2583_(_0125_, rst);
    not _2584_(_0126_, rst);
    not _2585_(_0127_, rst);
    not _2586_(_0128_, rst);
    not _2587_(_0129_, rst);
    not _2588_(_0130_, rst);
    not _2589_(_0131_, rst);
    not _2590_(_0132_, rst);
    not _2591_(_0133_, rst);
    not _2592_(_0134_, rst);
    not _2593_(_0135_, rst);
    not _2594_(_0136_, rst);
    not _2595_(_0137_, rst);
    not _2596_(_0138_, rst);
    not _2597_(_0139_, rst);
    not _2598_(_0140_, rst);
    not _2599_(_0141_, rst);
    not _2600_(_0142_, rst);
    not _2601_(_0143_, rst);
    not _2602_(_0144_, rst);
    not _2603_(_0145_, rst);
    not _2604_(_0146_, rst);
    not _2605_(_0147_, rst);
    not _2606_(_0148_, rst);
    not _2607_(_0149_, rst);
    not _2608_(_0150_, rst);
    not _2609_(_0151_, rst);
    not _2610_(_0152_, rst);
    not _2611_(_0153_, rst);
    not _2612_(_0154_, rst);
    not _2613_(_0155_, rst);
    not _2614_(_0156_, rst);
    not _2615_(_0157_, rst);
    not _2616_(_0158_, rst);
    not _2617_(_0159_, rst);
    not _2618_(_0160_, rst);
    not _2619_(_0161_, rst);
    not _2620_(_0162_, rst);
    not _2621_(_0163_, rst);
    not _2622_(_0164_, rst);
    not _2623_(_0165_, rst);
    not _2624_(_0166_, rst);
    not _2625_(_0167_, rst);
    not _2626_(_0168_, rst);
    not _2627_(_0169_, rst);
    not _2628_(_0170_, rst);
    not _2629_(_0171_, rst);
    not _2630_(_0172_, rst);
    not _2631_(_0173_, rst);
    not _2632_(_0174_, rst);
    not _2633_(_0175_, rst);
    not _2634_(_0176_, rst);
    not _2635_(_0177_, rst);
    not _2636_(_0178_, rst);
    not _2637_(_0179_, rst);
    not _2638_(_0180_, rst);
    not _2639_(_0181_, rst);
    not _2640_(_0182_, rst);
    not _2641_(_0183_, rst);
    not _2642_(_0184_, rst);
    not _2643_(_0185_, rst);
    not _2644_(_0186_, rst);
    not _2645_(_0187_, rst);
    not _2646_(_0188_, rst);
    not _2647_(_0189_, rst);
    not _2648_(_0190_, rst);
    dff _2649_(.RN(_0000_), .SN(1'b1), .CK(clk), .D(_0191_), .Q(\cache_tags[6][0]));
    dff _2650_(.RN(_0001_), .SN(1'b1), .CK(clk), .D(_0192_), .Q(\cache_tags[6][1]));
    dff _2651_(.RN(_0002_), .SN(1'b1), .CK(clk), .D(_0193_), .Q(\cache_tags[6][2]));
    dff _2652_(.RN(_0003_), .SN(1'b1), .CK(clk), .D(_0194_), .Q(\cache_tags[6][3]));
    dff _2653_(.RN(_0004_), .SN(1'b1), .CK(clk), .D(_0195_), .Q(cache_ready));
    dff _2654_(.RN(_0005_), .SN(1'b1), .CK(clk), .D(_0196_), .Q(cache_state[0]));
    dff _2655_(.RN(_0006_), .SN(1'b1), .CK(clk), .D(_0197_), .Q(cache_state[1]));
    dff _2656_(.RN(_0007_), .SN(1'b1), .CK(clk), .D(_0198_), .Q(cache_state[2]));
    dff _2657_(.RN(_0008_), .SN(1'b1), .CK(clk), .D(_0199_), .Q(access_index[0]));
    dff _2658_(.RN(_0009_), .SN(1'b1), .CK(clk), .D(_0200_), .Q(access_index[1]));
    dff _2659_(.RN(_0010_), .SN(1'b1), .CK(clk), .D(_0201_), .Q(access_index[2]));
    dff _2660_(.RN(_0011_), .SN(1'b1), .CK(clk), .D(_0202_), .Q(\cache_data[1][0]));
    dff _2661_(.RN(_0012_), .SN(1'b1), .CK(clk), .D(_0203_), .Q(\cache_data[1][1]));
    dff _2662_(.RN(_0013_), .SN(1'b1), .CK(clk), .D(_0204_), .Q(\cache_data[1][2]));
    dff _2663_(.RN(_0014_), .SN(1'b1), .CK(clk), .D(_0205_), .Q(\cache_data[1][3]));
    dff _2664_(.RN(_0015_), .SN(1'b1), .CK(clk), .D(_0206_), .Q(\cache_data[1][4]));
    dff _2665_(.RN(_0016_), .SN(1'b1), .CK(clk), .D(_0207_), .Q(\cache_data[1][5]));
    dff _2666_(.RN(_0017_), .SN(1'b1), .CK(clk), .D(_0208_), .Q(\cache_data[1][6]));
    dff _2667_(.RN(_0018_), .SN(1'b1), .CK(clk), .D(_0209_), .Q(\cache_data[1][7]));
    dff _2668_(.RN(_0019_), .SN(1'b1), .CK(clk), .D(_0210_), .Q(\cache_data[1][8]));
    dff _2669_(.RN(_0020_), .SN(1'b1), .CK(clk), .D(_0211_), .Q(\cache_data[1][9]));
    dff _2670_(.RN(_0021_), .SN(1'b1), .CK(clk), .D(_0212_), .Q(\cache_data[1][10]));
    dff _2671_(.RN(_0022_), .SN(1'b1), .CK(clk), .D(_0213_), .Q(\cache_data[1][11]));
    dff _2672_(.RN(_0023_), .SN(1'b1), .CK(clk), .D(_0214_), .Q(\cache_data[1][12]));
    dff _2673_(.RN(_0024_), .SN(1'b1), .CK(clk), .D(_0215_), .Q(\cache_data[1][13]));
    dff _2674_(.RN(_0025_), .SN(1'b1), .CK(clk), .D(_0216_), .Q(\cache_data[1][14]));
    dff _2675_(.RN(_0026_), .SN(1'b1), .CK(clk), .D(_0217_), .Q(\cache_data[1][15]));
    dff _2676_(.RN(_0027_), .SN(1'b1), .CK(clk), .D(_0218_), .Q(\cache_data[2][0]));
    dff _2677_(.RN(_0028_), .SN(1'b1), .CK(clk), .D(_0219_), .Q(\cache_data[2][1]));
    dff _2678_(.RN(_0029_), .SN(1'b1), .CK(clk), .D(_0220_), .Q(\cache_data[2][2]));
    dff _2679_(.RN(_0030_), .SN(1'b1), .CK(clk), .D(_0221_), .Q(\cache_data[2][3]));
    dff _2680_(.RN(_0031_), .SN(1'b1), .CK(clk), .D(_0222_), .Q(\cache_data[2][4]));
    dff _2681_(.RN(_0032_), .SN(1'b1), .CK(clk), .D(_0223_), .Q(\cache_data[2][5]));
    dff _2682_(.RN(_0033_), .SN(1'b1), .CK(clk), .D(_0224_), .Q(\cache_data[2][6]));
    dff _2683_(.RN(_0034_), .SN(1'b1), .CK(clk), .D(_0225_), .Q(\cache_data[2][7]));
    dff _2684_(.RN(_0035_), .SN(1'b1), .CK(clk), .D(_0226_), .Q(\cache_data[2][8]));
    dff _2685_(.RN(_0036_), .SN(1'b1), .CK(clk), .D(_0227_), .Q(\cache_data[2][9]));
    dff _2686_(.RN(_0037_), .SN(1'b1), .CK(clk), .D(_0228_), .Q(\cache_data[2][10]));
    dff _2687_(.RN(_0038_), .SN(1'b1), .CK(clk), .D(_0229_), .Q(\cache_data[2][11]));
    dff _2688_(.RN(_0039_), .SN(1'b1), .CK(clk), .D(_0230_), .Q(\cache_data[2][12]));
    dff _2689_(.RN(_0040_), .SN(1'b1), .CK(clk), .D(_0231_), .Q(\cache_data[2][13]));
    dff _2690_(.RN(_0041_), .SN(1'b1), .CK(clk), .D(_0232_), .Q(\cache_data[2][14]));
    dff _2691_(.RN(_0042_), .SN(1'b1), .CK(clk), .D(_0233_), .Q(\cache_data[2][15]));
    dff _2692_(.RN(_0043_), .SN(1'b1), .CK(clk), .D(_0234_), .Q(\cache_data[4][0]));
    dff _2693_(.RN(_0044_), .SN(1'b1), .CK(clk), .D(_0235_), .Q(\cache_data[4][1]));
    dff _2694_(.RN(_0045_), .SN(1'b1), .CK(clk), .D(_0236_), .Q(\cache_data[4][2]));
    dff _2695_(.RN(_0046_), .SN(1'b1), .CK(clk), .D(_0237_), .Q(\cache_data[4][3]));
    dff _2696_(.RN(_0047_), .SN(1'b1), .CK(clk), .D(_0238_), .Q(\cache_data[4][4]));
    dff _2697_(.RN(_0048_), .SN(1'b1), .CK(clk), .D(_0239_), .Q(\cache_data[4][5]));
    dff _2698_(.RN(_0049_), .SN(1'b1), .CK(clk), .D(_0240_), .Q(\cache_data[4][6]));
    dff _2699_(.RN(_0050_), .SN(1'b1), .CK(clk), .D(_0241_), .Q(\cache_data[4][7]));
    dff _2700_(.RN(_0051_), .SN(1'b1), .CK(clk), .D(_0242_), .Q(\cache_data[4][8]));
    dff _2701_(.RN(_0052_), .SN(1'b1), .CK(clk), .D(_0243_), .Q(\cache_data[4][9]));
    dff _2702_(.RN(_0053_), .SN(1'b1), .CK(clk), .D(_0244_), .Q(\cache_data[4][10]));
    dff _2703_(.RN(_0054_), .SN(1'b1), .CK(clk), .D(_0245_), .Q(\cache_data[4][11]));
    dff _2704_(.RN(_0055_), .SN(1'b1), .CK(clk), .D(_0246_), .Q(\cache_data[4][12]));
    dff _2705_(.RN(_0056_), .SN(1'b1), .CK(clk), .D(_0247_), .Q(\cache_data[4][13]));
    dff _2706_(.RN(_0057_), .SN(1'b1), .CK(clk), .D(_0248_), .Q(\cache_data[4][14]));
    dff _2707_(.RN(_0058_), .SN(1'b1), .CK(clk), .D(_0249_), .Q(\cache_data[4][15]));
    dff _2708_(.RN(_0059_), .SN(1'b1), .CK(clk), .D(_0250_), .Q(\cache_data[5][0]));
    dff _2709_(.RN(_0060_), .SN(1'b1), .CK(clk), .D(_0251_), .Q(\cache_data[5][1]));
    dff _2710_(.RN(_0061_), .SN(1'b1), .CK(clk), .D(_0252_), .Q(\cache_data[5][2]));
    dff _2711_(.RN(_0062_), .SN(1'b1), .CK(clk), .D(_0253_), .Q(\cache_data[5][3]));
    dff _2712_(.RN(_0063_), .SN(1'b1), .CK(clk), .D(_0254_), .Q(\cache_data[5][4]));
    dff _2713_(.RN(_0064_), .SN(1'b1), .CK(clk), .D(_0255_), .Q(\cache_data[5][5]));
    dff _2714_(.RN(_0065_), .SN(1'b1), .CK(clk), .D(_0256_), .Q(\cache_data[5][6]));
    dff _2715_(.RN(_0066_), .SN(1'b1), .CK(clk), .D(_0257_), .Q(\cache_data[5][7]));
    dff _2716_(.RN(_0067_), .SN(1'b1), .CK(clk), .D(_0258_), .Q(\cache_data[5][8]));
    dff _2717_(.RN(_0068_), .SN(1'b1), .CK(clk), .D(_0259_), .Q(\cache_data[5][9]));
    dff _2718_(.RN(_0069_), .SN(1'b1), .CK(clk), .D(_0260_), .Q(\cache_data[5][10]));
    dff _2719_(.RN(_0070_), .SN(1'b1), .CK(clk), .D(_0261_), .Q(\cache_data[5][11]));
    dff _2720_(.RN(_0071_), .SN(1'b1), .CK(clk), .D(_0262_), .Q(\cache_data[5][12]));
    dff _2721_(.RN(_0072_), .SN(1'b1), .CK(clk), .D(_0263_), .Q(\cache_data[5][13]));
    dff _2722_(.RN(_0073_), .SN(1'b1), .CK(clk), .D(_0264_), .Q(\cache_data[5][14]));
    dff _2723_(.RN(_0074_), .SN(1'b1), .CK(clk), .D(_0265_), .Q(\cache_data[5][15]));
    dff _2724_(.RN(_0075_), .SN(1'b1), .CK(clk), .D(_0266_), .Q(\cache_data[6][0]));
    dff _2725_(.RN(_0076_), .SN(1'b1), .CK(clk), .D(_0267_), .Q(\cache_data[6][1]));
    dff _2726_(.RN(_0077_), .SN(1'b1), .CK(clk), .D(_0268_), .Q(\cache_data[6][2]));
    dff _2727_(.RN(_0078_), .SN(1'b1), .CK(clk), .D(_0269_), .Q(\cache_data[6][3]));
    dff _2728_(.RN(_0079_), .SN(1'b1), .CK(clk), .D(_0270_), .Q(\cache_data[6][4]));
    dff _2729_(.RN(_0080_), .SN(1'b1), .CK(clk), .D(_0271_), .Q(\cache_data[6][5]));
    dff _2730_(.RN(_0081_), .SN(1'b1), .CK(clk), .D(_0272_), .Q(\cache_data[6][6]));
    dff _2731_(.RN(_0082_), .SN(1'b1), .CK(clk), .D(_0273_), .Q(\cache_data[6][7]));
    dff _2732_(.RN(_0083_), .SN(1'b1), .CK(clk), .D(_0274_), .Q(\cache_data[6][8]));
    dff _2733_(.RN(_0084_), .SN(1'b1), .CK(clk), .D(_0275_), .Q(\cache_data[6][9]));
    dff _2734_(.RN(_0085_), .SN(1'b1), .CK(clk), .D(_0276_), .Q(\cache_data[6][10]));
    dff _2735_(.RN(_0086_), .SN(1'b1), .CK(clk), .D(_0277_), .Q(\cache_data[6][11]));
    dff _2736_(.RN(_0087_), .SN(1'b1), .CK(clk), .D(_0278_), .Q(\cache_data[6][12]));
    dff _2737_(.RN(_0088_), .SN(1'b1), .CK(clk), .D(_0279_), .Q(\cache_data[6][13]));
    dff _2738_(.RN(_0089_), .SN(1'b1), .CK(clk), .D(_0280_), .Q(\cache_data[6][14]));
    dff _2739_(.RN(_0090_), .SN(1'b1), .CK(clk), .D(_0281_), .Q(\cache_data[6][15]));
    dff _2740_(.RN(_0091_), .SN(1'b1), .CK(clk), .D(_0282_), .Q(\cache_data[7][0]));
    dff _2741_(.RN(_0092_), .SN(1'b1), .CK(clk), .D(_0283_), .Q(\cache_data[7][1]));
    dff _2742_(.RN(_0093_), .SN(1'b1), .CK(clk), .D(_0284_), .Q(\cache_data[7][2]));
    dff _2743_(.RN(_0094_), .SN(1'b1), .CK(clk), .D(_0285_), .Q(\cache_data[7][3]));
    dff _2744_(.RN(_0095_), .SN(1'b1), .CK(clk), .D(_0286_), .Q(\cache_data[7][4]));
    dff _2745_(.RN(_0096_), .SN(1'b1), .CK(clk), .D(_0287_), .Q(\cache_data[7][5]));
    dff _2746_(.RN(_0097_), .SN(1'b1), .CK(clk), .D(_0288_), .Q(\cache_data[7][6]));
    dff _2747_(.RN(_0098_), .SN(1'b1), .CK(clk), .D(_0289_), .Q(\cache_data[7][7]));
    dff _2748_(.RN(_0099_), .SN(1'b1), .CK(clk), .D(_0290_), .Q(\cache_data[7][8]));
    dff _2749_(.RN(_0100_), .SN(1'b1), .CK(clk), .D(_0291_), .Q(\cache_data[7][9]));
    dff _2750_(.RN(_0101_), .SN(1'b1), .CK(clk), .D(_0292_), .Q(\cache_data[7][10]));
    dff _2751_(.RN(_0102_), .SN(1'b1), .CK(clk), .D(_0293_), .Q(\cache_data[7][11]));
    dff _2752_(.RN(_0103_), .SN(1'b1), .CK(clk), .D(_0294_), .Q(\cache_data[7][12]));
    dff _2753_(.RN(_0104_), .SN(1'b1), .CK(clk), .D(_0295_), .Q(\cache_data[7][13]));
    dff _2754_(.RN(_0105_), .SN(1'b1), .CK(clk), .D(_0296_), .Q(\cache_data[7][14]));
    dff _2755_(.RN(_0106_), .SN(1'b1), .CK(clk), .D(_0297_), .Q(\cache_data[7][15]));
    dff _2756_(.RN(_0107_), .SN(1'b1), .CK(clk), .D(_0298_), .Q(\cache_tags[0][0]));
    dff _2757_(.RN(_0108_), .SN(1'b1), .CK(clk), .D(_0299_), .Q(\cache_tags[0][1]));
    dff _2758_(.RN(_0109_), .SN(1'b1), .CK(clk), .D(_0300_), .Q(\cache_tags[0][2]));
    dff _2759_(.RN(_0110_), .SN(1'b1), .CK(clk), .D(_0301_), .Q(\cache_tags[0][3]));
    dff _2760_(.RN(_0111_), .SN(1'b1), .CK(clk), .D(_0302_), .Q(\cache_tags[1][0]));
    dff _2761_(.RN(_0112_), .SN(1'b1), .CK(clk), .D(_0303_), .Q(\cache_tags[1][1]));
    dff _2762_(.RN(_0113_), .SN(1'b1), .CK(clk), .D(_0304_), .Q(\cache_tags[1][2]));
    dff _2763_(.RN(_0114_), .SN(1'b1), .CK(clk), .D(_0305_), .Q(\cache_tags[1][3]));
    dff _2764_(.RN(_0115_), .SN(1'b1), .CK(clk), .D(_0306_), .Q(\cache_tags[2][0]));
    dff _2765_(.RN(_0116_), .SN(1'b1), .CK(clk), .D(_0307_), .Q(\cache_tags[2][1]));
    dff _2766_(.RN(_0117_), .SN(1'b1), .CK(clk), .D(_0308_), .Q(\cache_tags[2][2]));
    dff _2767_(.RN(_0118_), .SN(1'b1), .CK(clk), .D(_0309_), .Q(\cache_tags[2][3]));
    dff _2768_(.RN(_0119_), .SN(1'b1), .CK(clk), .D(_0310_), .Q(\cache_tags[3][0]));
    dff _2769_(.RN(_0120_), .SN(1'b1), .CK(clk), .D(_0311_), .Q(\cache_tags[3][1]));
    dff _2770_(.RN(_0121_), .SN(1'b1), .CK(clk), .D(_0312_), .Q(\cache_tags[3][2]));
    dff _2771_(.RN(_0122_), .SN(1'b1), .CK(clk), .D(_0313_), .Q(\cache_tags[3][3]));
    dff _2772_(.RN(_0123_), .SN(1'b1), .CK(clk), .D(_0314_), .Q(\cache_tags[4][0]));
    dff _2773_(.RN(_0124_), .SN(1'b1), .CK(clk), .D(_0315_), .Q(\cache_tags[4][1]));
    dff _2774_(.RN(_0125_), .SN(1'b1), .CK(clk), .D(_0316_), .Q(\cache_tags[4][2]));
    dff _2775_(.RN(_0126_), .SN(1'b1), .CK(clk), .D(_0317_), .Q(\cache_tags[4][3]));
    dff _2776_(.RN(_0127_), .SN(1'b1), .CK(clk), .D(_0318_), .Q(\cache_tags[5][0]));
    dff _2777_(.RN(_0128_), .SN(1'b1), .CK(clk), .D(_0319_), .Q(\cache_tags[5][1]));
    dff _2778_(.RN(_0129_), .SN(1'b1), .CK(clk), .D(_0320_), .Q(\cache_tags[5][2]));
    dff _2779_(.RN(_0130_), .SN(1'b1), .CK(clk), .D(_0321_), .Q(\cache_tags[5][3]));
    dff _2780_(.RN(_0131_), .SN(1'b1), .CK(clk), .D(_0322_), .Q(read_data[0]));
    dff _2781_(.RN(_0132_), .SN(1'b1), .CK(clk), .D(_0323_), .Q(read_data[1]));
    dff _2782_(.RN(_0133_), .SN(1'b1), .CK(clk), .D(_0324_), .Q(read_data[2]));
    dff _2783_(.RN(_0134_), .SN(1'b1), .CK(clk), .D(_0325_), .Q(read_data[3]));
    dff _2784_(.RN(_0135_), .SN(1'b1), .CK(clk), .D(_0326_), .Q(read_data[4]));
    dff _2785_(.RN(_0136_), .SN(1'b1), .CK(clk), .D(_0327_), .Q(read_data[5]));
    dff _2786_(.RN(_0137_), .SN(1'b1), .CK(clk), .D(_0328_), .Q(read_data[6]));
    dff _2787_(.RN(_0138_), .SN(1'b1), .CK(clk), .D(_0329_), .Q(read_data[7]));
    dff _2788_(.RN(_0139_), .SN(1'b1), .CK(clk), .D(_0330_), .Q(read_data[8]));
    dff _2789_(.RN(_0140_), .SN(1'b1), .CK(clk), .D(_0331_), .Q(read_data[9]));
    dff _2790_(.RN(_0141_), .SN(1'b1), .CK(clk), .D(_0332_), .Q(read_data[10]));
    dff _2791_(.RN(_0142_), .SN(1'b1), .CK(clk), .D(_0333_), .Q(read_data[11]));
    dff _2792_(.RN(_0143_), .SN(1'b1), .CK(clk), .D(_0334_), .Q(read_data[12]));
    dff _2793_(.RN(_0144_), .SN(1'b1), .CK(clk), .D(_0335_), .Q(read_data[13]));
    dff _2794_(.RN(_0145_), .SN(1'b1), .CK(clk), .D(_0336_), .Q(read_data[14]));
    dff _2795_(.RN(_0146_), .SN(1'b1), .CK(clk), .D(_0337_), .Q(read_data[15]));
    dff _2796_(.RN(_0147_), .SN(1'b1), .CK(clk), .D(_0338_), .Q(\cache_tags[7][0]));
    dff _2797_(.RN(_0148_), .SN(1'b1), .CK(clk), .D(_0339_), .Q(\cache_tags[7][1]));
    dff _2798_(.RN(_0149_), .SN(1'b1), .CK(clk), .D(_0340_), .Q(\cache_tags[7][2]));
    dff _2799_(.RN(_0150_), .SN(1'b1), .CK(clk), .D(_0341_), .Q(\cache_tags[7][3]));
    dff _2800_(.RN(_0151_), .SN(1'b1), .CK(clk), .D(_0342_), .Q(\cache_data[3][0]));
    dff _2801_(.RN(_0152_), .SN(1'b1), .CK(clk), .D(_0343_), .Q(\cache_data[3][1]));
    dff _2802_(.RN(_0153_), .SN(1'b1), .CK(clk), .D(_0344_), .Q(\cache_data[3][2]));
    dff _2803_(.RN(_0154_), .SN(1'b1), .CK(clk), .D(_0345_), .Q(\cache_data[3][3]));
    dff _2804_(.RN(_0155_), .SN(1'b1), .CK(clk), .D(_0346_), .Q(\cache_data[3][4]));
    dff _2805_(.RN(_0156_), .SN(1'b1), .CK(clk), .D(_0347_), .Q(\cache_data[3][5]));
    dff _2806_(.RN(_0157_), .SN(1'b1), .CK(clk), .D(_0348_), .Q(\cache_data[3][6]));
    dff _2807_(.RN(_0158_), .SN(1'b1), .CK(clk), .D(_0349_), .Q(\cache_data[3][7]));
    dff _2808_(.RN(_0159_), .SN(1'b1), .CK(clk), .D(_0350_), .Q(\cache_data[3][8]));
    dff _2809_(.RN(_0160_), .SN(1'b1), .CK(clk), .D(_0351_), .Q(\cache_data[3][9]));
    dff _2810_(.RN(_0161_), .SN(1'b1), .CK(clk), .D(_0352_), .Q(\cache_data[3][10]));
    dff _2811_(.RN(_0162_), .SN(1'b1), .CK(clk), .D(_0353_), .Q(\cache_data[3][11]));
    dff _2812_(.RN(_0163_), .SN(1'b1), .CK(clk), .D(_0354_), .Q(\cache_data[3][12]));
    dff _2813_(.RN(_0164_), .SN(1'b1), .CK(clk), .D(_0355_), .Q(\cache_data[3][13]));
    dff _2814_(.RN(_0165_), .SN(1'b1), .CK(clk), .D(_0356_), .Q(\cache_data[3][14]));
    dff _2815_(.RN(_0166_), .SN(1'b1), .CK(clk), .D(_0357_), .Q(\cache_data[3][15]));
    dff _2816_(.RN(_0167_), .SN(1'b1), .CK(clk), .D(_0358_), .Q(\cache_data[0][0]));
    dff _2817_(.RN(_0168_), .SN(1'b1), .CK(clk), .D(_0359_), .Q(\cache_data[0][1]));
    dff _2818_(.RN(_0169_), .SN(1'b1), .CK(clk), .D(_0360_), .Q(\cache_data[0][2]));
    dff _2819_(.RN(_0170_), .SN(1'b1), .CK(clk), .D(_0361_), .Q(\cache_data[0][3]));
    dff _2820_(.RN(_0171_), .SN(1'b1), .CK(clk), .D(_0362_), .Q(\cache_data[0][4]));
    dff _2821_(.RN(_0172_), .SN(1'b1), .CK(clk), .D(_0363_), .Q(\cache_data[0][5]));
    dff _2822_(.RN(_0173_), .SN(1'b1), .CK(clk), .D(_0364_), .Q(\cache_data[0][6]));
    dff _2823_(.RN(_0174_), .SN(1'b1), .CK(clk), .D(_0365_), .Q(\cache_data[0][7]));
    dff _2824_(.RN(_0175_), .SN(1'b1), .CK(clk), .D(_0366_), .Q(\cache_data[0][8]));
    dff _2825_(.RN(_0176_), .SN(1'b1), .CK(clk), .D(_0367_), .Q(\cache_data[0][9]));
    dff _2826_(.RN(_0177_), .SN(1'b1), .CK(clk), .D(_0368_), .Q(\cache_data[0][10]));
    dff _2827_(.RN(_0178_), .SN(1'b1), .CK(clk), .D(_0369_), .Q(\cache_data[0][11]));
    dff _2828_(.RN(_0179_), .SN(1'b1), .CK(clk), .D(_0370_), .Q(\cache_data[0][12]));
    dff _2829_(.RN(_0180_), .SN(1'b1), .CK(clk), .D(_0371_), .Q(\cache_data[0][13]));
    dff _2830_(.RN(_0181_), .SN(1'b1), .CK(clk), .D(_0372_), .Q(\cache_data[0][14]));
    dff _2831_(.RN(_0182_), .SN(1'b1), .CK(clk), .D(_0373_), .Q(\cache_data[0][15]));
    dff _2832_(.RN(_0183_), .SN(1'b1), .CK(clk), .D(_0374_), .Q(valid_bits[0]));
    dff _2833_(.RN(_0184_), .SN(1'b1), .CK(clk), .D(_0375_), .Q(valid_bits[1]));
    dff _2834_(.RN(_0185_), .SN(1'b1), .CK(clk), .D(_0376_), .Q(valid_bits[2]));
    dff _2835_(.RN(_0186_), .SN(1'b1), .CK(clk), .D(_0377_), .Q(valid_bits[3]));
    dff _2836_(.RN(_0187_), .SN(1'b1), .CK(clk), .D(_0378_), .Q(valid_bits[4]));
    dff _2837_(.RN(_0188_), .SN(1'b1), .CK(clk), .D(_0379_), .Q(valid_bits[5]));
    dff _2838_(.RN(_0189_), .SN(1'b1), .CK(clk), .D(_0380_), .Q(valid_bits[6]));
    dff _2839_(.RN(_0190_), .SN(1'b1), .CK(clk), .D(_0381_), .Q(valid_bits[7]));
endmodule