module trojan0_counter_host_0001(clk, rst, enable, count_out, overflow, pulse_out);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  wire _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire _142_;
  wire _143_;
  wire _144_;
  wire _145_;
  wire _146_;
  wire _147_;
  wire _148_;
  wire _149_;
  wire _150_;
  wire _151_;
  wire _152_;
  wire _153_;
  wire _154_;
  wire _155_;
  wire _156_;
  wire _157_;
  wire _158_;
  wire _159_;
  wire _160_;
  wire _161_;
  wire _162_;
  wire _163_;
  wire _164_;
  wire _165_;
  wire _166_;
  wire _167_;
  wire _168_;
  wire _169_;
  wire _170_;
  wire _171_;
  wire _172_;
  wire _173_;
  wire _174_;
  wire _175_;
  wire _176_;
  wire _177_;
  wire _178_;
  wire _179_;
  wire _180_;
  wire _181_;
  wire _182_;
  wire _183_;
  wire _184_;
  wire _185_;
  wire _186_;
  wire _187_;
  wire _188_;
  wire _189_;
  wire _190_;
  wire _191_;
  wire _192_;
  wire _193_;
  wire _194_;
  wire _195_;
  wire _196_;
  wire _197_;
  wire _198_;
  wire _199_;
  wire _200_;
  wire _201_;
  wire _202_;
  wire _203_;
  wire _204_;
  wire _205_;
  wire _206_;
  wire _207_;
  wire _208_;
  input clk;
  wire clk;
  output [11:0] count_out;
  wire [11:0] count_out;
  wire [11:0] counter;
  input enable;
  wire enable;
  output overflow;
  wire overflow;
  wire [11:0] period_counter;
  output pulse_out;
  wire pulse_out;
  input rst;
  wire rst;
    not _209_(_000_, rst);
    not _210_(_203_, enable);
    and _211_(_204_, _203_, overflow);
    and _212_(_205_, counter[1], counter[0]);
    and _213_(_206_, counter[3], counter[2]);
    and _214_(_207_, _206_, _205_);
    and _215_(_208_, counter[5], counter[4]);
    and _216_(_064_, counter[7], counter[6]);
    and _217_(_065_, _064_, _208_);
    and _218_(_066_, _065_, _207_);
    and _219_(_067_, counter[9], counter[8]);
    and _220_(_068_, counter[11], counter[10]);
    and _221_(_069_, _068_, _067_);
    and _222_(_070_, _069_, _066_);
    and _223_(_071_, _070_, enable);
    or _224_(_038_, _071_, _204_);
    and _225_(_072_, pulse_out, _203_);
    nor _226_(_073_, period_counter[11], period_counter[10]);
    nor _227_(_074_, period_counter[9], period_counter[8]);
    and _228_(_075_, _074_, _073_);
    not _229_(_076_, period_counter[7]);
    and _230_(_077_, _076_, period_counter[6]);
    not _231_(_078_, period_counter[4]);
    and _232_(_079_, period_counter[5], _078_);
    and _233_(_080_, _079_, _077_);
    and _234_(_081_, period_counter[1], period_counter[0]);
    nor _235_(_082_, period_counter[3], period_counter[2]);
    nand _236_(_083_, _082_, _081_);
    not _237_(_084_, _083_);
    and _238_(_085_, _084_, _080_);
    nand _239_(_086_, _085_, _075_);
    nor _240_(_087_, period_counter[11], period_counter[10]);
    or _241_(_088_, period_counter[9], period_counter[8]);
    nand _242_(_089_, _088_, _073_);
    and _243_(_090_, _089_, _087_);
    and _244_(_091_, period_counter[5], period_counter[4]);
    nand _245_(_092_, _091_, _077_);
    and _246_(_093_, _092_, _076_);
    nor _247_(_094_, period_counter[3], period_counter[2]);
    nand _248_(_095_, _094_, _083_);
    nand _249_(_096_, _095_, _080_);
    nand _250_(_097_, _096_, _093_);
    nand _251_(_098_, _097_, _075_);
    and _252_(_099_, _098_, _090_);
    and _253_(_100_, _099_, _086_);
    nor _254_(_101_, _100_, _203_);
    or _255_(_039_, _101_, _072_);
    xor _256_(_040_, counter[0], enable);
    and _257_(_102_, counter[1], _203_);
    xor _258_(_103_, counter[1], counter[0]);
    and _259_(_104_, _103_, enable);
    or _260_(_041_, _104_, _102_);
    and _261_(_105_, counter[2], _203_);
    xor _262_(_106_, _205_, counter[2]);
    and _263_(_107_, _106_, enable);
    or _264_(_042_, _107_, _105_);
    and _265_(_108_, counter[3], _203_);
    and _266_(_109_, _205_, counter[2]);
    xor _267_(_110_, _109_, counter[3]);
    and _268_(_111_, _110_, enable);
    or _269_(_043_, _111_, _108_);
    and _270_(_112_, counter[4], _203_);
    xor _271_(_113_, _207_, counter[4]);
    and _272_(_114_, _113_, enable);
    or _273_(_044_, _114_, _112_);
    and _274_(_115_, counter[5], _203_);
    and _275_(_116_, _207_, counter[4]);
    xor _276_(_117_, _116_, counter[5]);
    and _277_(_118_, _117_, enable);
    or _278_(_045_, _118_, _115_);
    and _279_(_119_, counter[6], _203_);
    and _280_(_120_, _208_, _207_);
    xor _281_(_121_, _120_, counter[6]);
    and _282_(_122_, _121_, enable);
    or _283_(_046_, _122_, _119_);
    and _284_(_123_, counter[7], _203_);
    and _285_(_124_, _120_, counter[6]);
    xor _286_(_125_, _124_, counter[7]);
    and _287_(_126_, _125_, enable);
    or _288_(_047_, _126_, _123_);
    and _289_(_127_, counter[8], _203_);
    xor _290_(_128_, _066_, counter[8]);
    and _291_(_129_, _128_, enable);
    or _292_(_048_, _129_, _127_);
    and _293_(_130_, counter[9], _203_);
    and _294_(_131_, _066_, counter[8]);
    xor _295_(_132_, _131_, counter[9]);
    and _296_(_133_, _132_, enable);
    or _297_(_049_, _133_, _130_);
    and _298_(_134_, counter[10], _203_);
    and _299_(_135_, _067_, _066_);
    xor _300_(_136_, _135_, counter[10]);
    and _301_(_137_, _136_, enable);
    or _302_(_050_, _137_, _134_);
    and _303_(_138_, counter[11], _203_);
    and _304_(_139_, _135_, counter[10]);
    xor _305_(_140_, _139_, counter[11]);
    and _306_(_141_, _140_, enable);
    or _307_(_051_, _141_, _138_);
    and _308_(_142_, period_counter[0], _203_);
    not _309_(_143_, period_counter[0]);
    and _310_(_144_, _100_, _143_);
    and _311_(_145_, _144_, enable);
    or _312_(_052_, _145_, _142_);
    and _313_(_146_, period_counter[1], _203_);
    xor _314_(_147_, period_counter[1], period_counter[0]);
    and _315_(_148_, _147_, _100_);
    and _316_(_149_, _148_, enable);
    or _317_(_053_, _149_, _146_);
    and _318_(_150_, period_counter[2], _203_);
    xor _319_(_151_, _081_, period_counter[2]);
    and _320_(_152_, _151_, _100_);
    and _321_(_153_, _152_, enable);
    or _322_(_054_, _153_, _150_);
    and _323_(_154_, period_counter[3], _203_);
    and _324_(_155_, _081_, period_counter[2]);
    xor _325_(_156_, _155_, period_counter[3]);
    and _326_(_157_, _156_, _100_);
    and _327_(_158_, _157_, enable);
    or _328_(_055_, _158_, _154_);
    and _329_(_159_, period_counter[4], _203_);
    and _330_(_160_, period_counter[3], period_counter[2]);
    and _331_(_161_, _160_, _081_);
    xor _332_(_162_, _161_, period_counter[4]);
    and _333_(_163_, _162_, _100_);
    and _334_(_164_, _163_, enable);
    or _335_(_056_, _164_, _159_);
    and _336_(_165_, period_counter[5], _203_);
    and _337_(_166_, _161_, period_counter[4]);
    xor _338_(_167_, _166_, period_counter[5]);
    and _339_(_168_, _167_, _100_);
    and _340_(_169_, _168_, enable);
    or _341_(_057_, _169_, _165_);
    and _342_(_170_, period_counter[6], _203_);
    and _343_(_171_, _161_, _091_);
    xor _344_(_172_, _171_, period_counter[6]);
    and _345_(_173_, _172_, _100_);
    and _346_(_174_, _173_, enable);
    or _347_(_058_, _174_, _170_);
    and _348_(_175_, period_counter[7], _203_);
    and _349_(_176_, _171_, period_counter[6]);
    xor _350_(_177_, _176_, period_counter[7]);
    and _351_(_178_, _177_, _100_);
    and _352_(_179_, _178_, enable);
    or _353_(_059_, _179_, _175_);
    and _354_(_180_, period_counter[8], _203_);
    and _355_(_181_, period_counter[7], period_counter[6]);
    and _356_(_182_, _181_, _091_);
    and _357_(_183_, _182_, _161_);
    xor _358_(_184_, _183_, period_counter[8]);
    and _359_(_185_, _184_, _100_);
    and _360_(_186_, _185_, enable);
    or _361_(_060_, _186_, _180_);
    and _362_(_187_, period_counter[9], _203_);
    and _363_(_188_, _183_, period_counter[8]);
    xor _364_(_189_, _188_, period_counter[9]);
    and _365_(_190_, _189_, _100_);
    and _366_(_191_, _190_, enable);
    or _367_(_061_, _191_, _187_);
    and _368_(_192_, period_counter[10], _203_);
    and _369_(_193_, period_counter[9], period_counter[8]);
    and _370_(_194_, _193_, _183_);
    xor _371_(_195_, _194_, period_counter[10]);
    and _372_(_196_, _195_, _100_);
    and _373_(_197_, _196_, enable);
    or _374_(_062_, _197_, _192_);
    and _375_(_198_, period_counter[11], _203_);
    and _376_(_199_, _194_, period_counter[10]);
    xor _377_(_200_, _199_, period_counter[11]);
    and _378_(_201_, _200_, _100_);
    and _379_(_202_, _201_, enable);
    or _380_(_063_, _202_, _198_);
    not _381_(_001_, rst);
    not _382_(_002_, rst);
    not _383_(_003_, rst);
    not _384_(_004_, rst);
    not _385_(_005_, rst);
    not _386_(_006_, rst);
    not _387_(_007_, rst);
    not _388_(_008_, rst);
    not _389_(_009_, rst);
    not _390_(_010_, rst);
    not _391_(_011_, rst);
    not _392_(_012_, rst);
    not _393_(_013_, rst);
    not _394_(_014_, rst);
    not _395_(_015_, rst);
    not _396_(_016_, rst);
    not _397_(_017_, rst);
    not _398_(_018_, rst);
    not _399_(_019_, rst);
    not _400_(_020_, rst);
    not _401_(_021_, rst);
    not _402_(_022_, rst);
    not _403_(_023_, rst);
    not _404_(_024_, rst);
    not _405_(_025_, rst);
    not _406_(_026_, rst);
    not _407_(_027_, rst);
    not _408_(_028_, rst);
    not _409_(_029_, rst);
    not _410_(_030_, rst);
    not _411_(_031_, rst);
    not _412_(_032_, rst);
    not _413_(_033_, rst);
    not _414_(_034_, rst);
    not _415_(_035_, rst);
    not _416_(_036_, rst);
    not _417_(_037_, rst);
    dff _418_(.RN(_000_), .SN(1'b1), .CK(clk), .D(_038_), .Q(overflow));
    dff _419_(.RN(_001_), .SN(1'b1), .CK(clk), .D(counter[0]), .Q(count_out[0]));
    dff _420_(.RN(_002_), .SN(1'b1), .CK(clk), .D(counter[1]), .Q(count_out[1]));
    dff _421_(.RN(_003_), .SN(1'b1), .CK(clk), .D(counter[2]), .Q(count_out[2]));
    dff _422_(.RN(_004_), .SN(1'b1), .CK(clk), .D(counter[3]), .Q(count_out[3]));
    dff _423_(.RN(_005_), .SN(1'b1), .CK(clk), .D(counter[4]), .Q(count_out[4]));
    dff _424_(.RN(_006_), .SN(1'b1), .CK(clk), .D(counter[5]), .Q(count_out[5]));
    dff _425_(.RN(_007_), .SN(1'b1), .CK(clk), .D(counter[6]), .Q(count_out[6]));
    dff _426_(.RN(_008_), .SN(1'b1), .CK(clk), .D(counter[7]), .Q(count_out[7]));
    dff _427_(.RN(_009_), .SN(1'b1), .CK(clk), .D(counter[8]), .Q(count_out[8]));
    dff _428_(.RN(_010_), .SN(1'b1), .CK(clk), .D(counter[9]), .Q(count_out[9]));
    dff _429_(.RN(_011_), .SN(1'b1), .CK(clk), .D(counter[10]), .Q(count_out[10]));
    dff _430_(.RN(_012_), .SN(1'b1), .CK(clk), .D(counter[11]), .Q(count_out[11]));
    dff _431_(.RN(_013_), .SN(1'b1), .CK(clk), .D(_039_), .Q(pulse_out));
    dff _432_(.RN(_014_), .SN(1'b1), .CK(clk), .D(_040_), .Q(counter[0]));
    dff _433_(.RN(_015_), .SN(1'b1), .CK(clk), .D(_041_), .Q(counter[1]));
    dff _434_(.RN(_016_), .SN(1'b1), .CK(clk), .D(_042_), .Q(counter[2]));
    dff _435_(.RN(_017_), .SN(1'b1), .CK(clk), .D(_043_), .Q(counter[3]));
    dff _436_(.RN(_018_), .SN(1'b1), .CK(clk), .D(_044_), .Q(counter[4]));
    dff _437_(.RN(_019_), .SN(1'b1), .CK(clk), .D(_045_), .Q(counter[5]));
    dff _438_(.RN(_020_), .SN(1'b1), .CK(clk), .D(_046_), .Q(counter[6]));
    dff _439_(.RN(_021_), .SN(1'b1), .CK(clk), .D(_047_), .Q(counter[7]));
    dff _440_(.RN(_022_), .SN(1'b1), .CK(clk), .D(_048_), .Q(counter[8]));
    dff _441_(.RN(_023_), .SN(1'b1), .CK(clk), .D(_049_), .Q(counter[9]));
    dff _442_(.RN(_024_), .SN(1'b1), .CK(clk), .D(_050_), .Q(counter[10]));
    dff _443_(.RN(_025_), .SN(1'b1), .CK(clk), .D(_051_), .Q(counter[11]));
    dff _444_(.RN(_026_), .SN(1'b1), .CK(clk), .D(_052_), .Q(period_counter[0]));
    dff _445_(.RN(_027_), .SN(1'b1), .CK(clk), .D(_053_), .Q(period_counter[1]));
    dff _446_(.RN(_028_), .SN(1'b1), .CK(clk), .D(_054_), .Q(period_counter[2]));
    dff _447_(.RN(_029_), .SN(1'b1), .CK(clk), .D(_055_), .Q(period_counter[3]));
    dff _448_(.RN(_030_), .SN(1'b1), .CK(clk), .D(_056_), .Q(period_counter[4]));
    dff _449_(.RN(_031_), .SN(1'b1), .CK(clk), .D(_057_), .Q(period_counter[5]));
    dff _450_(.RN(_032_), .SN(1'b1), .CK(clk), .D(_058_), .Q(period_counter[6]));
    dff _451_(.RN(_033_), .SN(1'b1), .CK(clk), .D(_059_), .Q(period_counter[7]));
    dff _452_(.RN(_034_), .SN(1'b1), .CK(clk), .D(_060_), .Q(period_counter[8]));
    dff _453_(.RN(_035_), .SN(1'b1), .CK(clk), .D(_061_), .Q(period_counter[9]));
    dff _454_(.RN(_036_), .SN(1'b1), .CK(clk), .D(_062_), .Q(period_counter[10]));
    dff _455_(.RN(_037_), .SN(1'b1), .CK(clk), .D(_063_), .Q(period_counter[11]));
endmodule