module trojan0_network_host_0001(clk, rst, packet_in, packet_valid, dest_addr, packet_out, packet_ready, route_error);
  wire _0000_;
  wire _0001_;
  wire _0002_;
  wire _0003_;
  wire _0004_;
  wire _0005_;
  wire _0006_;
  wire _0007_;
  wire _0008_;
  wire _0009_;
  wire _0010_;
  wire _0011_;
  wire _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  wire _0514_;
  wire _0515_;
  wire _0516_;
  wire _0517_;
  wire _0518_;
  wire _0519_;
  wire _0520_;
  wire _0521_;
  wire _0522_;
  wire _0523_;
  wire _0524_;
  wire _0525_;
  wire _0526_;
  wire _0527_;
  wire _0528_;
  wire _0529_;
  wire _0530_;
  wire _0531_;
  wire _0532_;
  wire _0533_;
  wire _0534_;
  wire _0535_;
  wire _0536_;
  wire _0537_;
  wire _0538_;
  wire _0539_;
  wire _0540_;
  wire _0541_;
  wire _0542_;
  wire _0543_;
  wire _0544_;
  wire _0545_;
  wire _0546_;
  wire _0547_;
  wire _0548_;
  wire _0549_;
  wire _0550_;
  wire _0551_;
  wire _0552_;
  wire _0553_;
  wire _0554_;
  wire _0555_;
  wire _0556_;
  wire _0557_;
  wire _0558_;
  wire _0559_;
  wire _0560_;
  wire _0561_;
  wire _0562_;
  wire _0563_;
  wire _0564_;
  wire _0565_;
  wire _0566_;
  wire _0567_;
  wire _0568_;
  wire _0569_;
  wire _0570_;
  wire _0571_;
  wire _0572_;
  wire _0573_;
  wire _0574_;
  wire _0575_;
  wire _0576_;
  wire _0577_;
  wire _0578_;
  wire _0579_;
  wire _0580_;
  wire _0581_;
  wire _0582_;
  wire _0583_;
  wire _0584_;
  wire _0585_;
  wire _0586_;
  wire _0587_;
  wire _0588_;
  wire _0589_;
  wire _0590_;
  wire _0591_;
  wire _0592_;
  wire _0593_;
  wire _0594_;
  wire _0595_;
  wire _0596_;
  wire _0597_;
  wire _0598_;
  wire _0599_;
  wire _0600_;
  wire _0601_;
  wire _0602_;
  wire _0603_;
  wire _0604_;
  wire _0605_;
  wire _0606_;
  wire _0607_;
  wire _0608_;
  wire _0609_;
  wire _0610_;
  wire _0611_;
  wire _0612_;
  wire _0613_;
  wire _0614_;
  wire _0615_;
  wire _0616_;
  wire _0617_;
  wire _0618_;
  wire _0619_;
  wire _0620_;
  wire _0621_;
  wire _0622_;
  wire _0623_;
  wire _0624_;
  wire _0625_;
  wire _0626_;
  wire _0627_;
  wire _0628_;
  wire _0629_;
  wire _0630_;
  wire _0631_;
  wire _0632_;
  wire _0633_;
  wire _0634_;
  wire _0635_;
  wire _0636_;
  wire _0637_;
  wire _0638_;
  wire _0639_;
  wire _0640_;
  wire _0641_;
  wire _0642_;
  wire _0643_;
  wire _0644_;
  wire _0645_;
  wire _0646_;
  wire _0647_;
  wire _0648_;
  wire _0649_;
  wire _0650_;
  wire _0651_;
  wire _0652_;
  wire _0653_;
  wire _0654_;
  wire _0655_;
  wire _0656_;
  wire _0657_;
  wire _0658_;
  wire _0659_;
  wire _0660_;
  wire _0661_;
  wire _0662_;
  wire _0663_;
  wire _0664_;
  wire _0665_;
  wire _0666_;
  wire _0667_;
  wire _0668_;
  wire _0669_;
  wire _0670_;
  wire _0671_;
  wire _0672_;
  wire _0673_;
  wire _0674_;
  wire _0675_;
  wire _0676_;
  wire _0677_;
  wire _0678_;
  wire _0679_;
  wire _0680_;
  wire _0681_;
  wire _0682_;
  wire _0683_;
  wire _0684_;
  wire _0685_;
  wire _0686_;
  wire _0687_;
  wire _0688_;
  wire _0689_;
  wire _0690_;
  wire _0691_;
  wire _0692_;
  wire _0693_;
  wire _0694_;
  wire _0695_;
  wire _0696_;
  wire _0697_;
  wire _0698_;
  wire _0699_;
  wire _0700_;
  wire _0701_;
  wire _0702_;
  wire _0703_;
  wire _0704_;
  wire _0705_;
  wire _0706_;
  wire _0707_;
  wire _0708_;
  wire _0709_;
  wire _0710_;
  wire _0711_;
  wire _0712_;
  wire _0713_;
  wire _0714_;
  wire _0715_;
  wire _0716_;
  wire _0717_;
  wire _0718_;
  wire _0719_;
  wire _0720_;
  wire _0721_;
  wire _0722_;
  wire _0723_;
  wire _0724_;
  wire _0725_;
  wire _0726_;
  wire _0727_;
  wire _0728_;
  wire _0729_;
  wire _0730_;
  wire _0731_;
  wire _0732_;
  wire _0733_;
  wire _0734_;
  wire _0735_;
  wire _0736_;
  wire _0737_;
  wire _0738_;
  wire _0739_;
  wire _0740_;
  wire _0741_;
  wire _0742_;
  wire _0743_;
  wire _0744_;
  wire _0745_;
  wire _0746_;
  wire _0747_;
  wire _0748_;
  wire _0749_;
  wire _0750_;
  wire _0751_;
  wire _0752_;
  wire _0753_;
  wire _0754_;
  wire _0755_;
  wire _0756_;
  wire _0757_;
  wire _0758_;
  wire _0759_;
  wire _0760_;
  wire _0761_;
  wire _0762_;
  wire _0763_;
  wire _0764_;
  wire _0765_;
  wire _0766_;
  wire _0767_;
  wire _0768_;
  wire _0769_;
  wire _0770_;
  wire _0771_;
  wire _0772_;
  wire _0773_;
  wire _0774_;
  wire _0775_;
  wire _0776_;
  wire _0777_;
  wire _0778_;
  wire _0779_;
  wire _0780_;
  wire _0781_;
  wire _0782_;
  wire _0783_;
  wire _0784_;
  wire _0785_;
  wire _0786_;
  wire _0787_;
  wire _0788_;
  wire _0789_;
  wire _0790_;
  wire _0791_;
  wire _0792_;
  wire _0793_;
  wire _0794_;
  wire _0795_;
  wire _0796_;
  wire _0797_;
  wire _0798_;
  wire _0799_;
  wire _0800_;
  wire _0801_;
  wire _0802_;
  wire _0803_;
  wire _0804_;
  wire _0805_;
  wire _0806_;
  wire _0807_;
  wire _0808_;
  wire _0809_;
  wire _0810_;
  wire _0811_;
  wire _0812_;
  wire _0813_;
  wire _0814_;
  wire _0815_;
  wire _0816_;
  wire _0817_;
  wire _0818_;
  wire _0819_;
  wire _0820_;
  wire _0821_;
  wire _0822_;
  wire _0823_;
  wire _0824_;
  wire _0825_;
  wire _0826_;
  wire _0827_;
  wire _0828_;
  wire _0829_;
  wire _0830_;
  wire _0831_;
  wire _0832_;
  wire _0833_;
  wire _0834_;
  wire _0835_;
  wire _0836_;
  wire _0837_;
  wire _0838_;
  wire _0839_;
  wire _0840_;
  wire _0841_;
  wire _0842_;
  wire _0843_;
  wire _0844_;
  wire _0845_;
  wire _0846_;
  wire _0847_;
  wire _0848_;
  wire _0849_;
  wire _0850_;
  wire _0851_;
  wire _0852_;
  wire _0853_;
  wire _0854_;
  wire _0855_;
  wire _0856_;
  wire _0857_;
  wire _0858_;
  wire _0859_;
  wire _0860_;
  wire _0861_;
  wire _0862_;
  wire _0863_;
  wire _0864_;
  wire _0865_;
  wire _0866_;
  wire _0867_;
  wire _0868_;
  wire _0869_;
  wire _0870_;
  wire _0871_;
  wire _0872_;
  wire _0873_;
  wire _0874_;
  wire _0875_;
  wire _0876_;
  wire _0877_;
  wire _0878_;
  wire _0879_;
  wire _0880_;
  wire _0881_;
  wire _0882_;
  wire _0883_;
  wire _0884_;
  wire _0885_;
  wire _0886_;
  wire _0887_;
  wire _0888_;
  wire _0889_;
  wire _0890_;
  wire _0891_;
  wire _0892_;
  wire _0893_;
  wire _0894_;
  wire _0895_;
  wire _0896_;
  wire _0897_;
  wire _0898_;
  wire _0899_;
  wire _0900_;
  wire _0901_;
  wire _0902_;
  wire _0903_;
  wire _0904_;
  wire _0905_;
  wire _0906_;
  wire _0907_;
  wire _0908_;
  wire _0909_;
  wire _0910_;
  wire _0911_;
  wire _0912_;
  wire _0913_;
  wire _0914_;
  wire _0915_;
  wire _0916_;
  wire _0917_;
  wire _0918_;
  wire _0919_;
  wire _0920_;
  wire _0921_;
  wire _0922_;
  wire _0923_;
  wire _0924_;
  wire _0925_;
  wire _0926_;
  wire _0927_;
  wire _0928_;
  wire _0929_;
  wire _0930_;
  wire _0931_;
  wire _0932_;
  wire _0933_;
  wire _0934_;
  wire _0935_;
  wire _0936_;
  wire _0937_;
  wire _0938_;
  wire _0939_;
  wire _0940_;
  wire _0941_;
  wire _0942_;
  wire _0943_;
  wire _0944_;
  wire _0945_;
  wire _0946_;
  wire _0947_;
  wire _0948_;
  wire _0949_;
  wire _0950_;
  wire _0951_;
  wire _0952_;
  wire _0953_;
  wire _0954_;
  wire _0955_;
  wire _0956_;
  wire _0957_;
  wire _0958_;
  wire _0959_;
  wire _0960_;
  wire _0961_;
  wire _0962_;
  wire _0963_;
  wire _0964_;
  wire _0965_;
  wire _0966_;
  wire _0967_;
  wire _0968_;
  wire _0969_;
  wire _0970_;
  wire _0971_;
  wire _0972_;
  wire _0973_;
  wire _0974_;
  wire _0975_;
  wire _0976_;
  wire _0977_;
  wire _0978_;
  wire _0979_;
  wire _0980_;
  wire _0981_;
  wire _0982_;
  wire _0983_;
  wire _0984_;
  wire _0985_;
  wire _0986_;
  wire _0987_;
  wire _0988_;
  wire _0989_;
  wire _0990_;
  wire _0991_;
  wire _0992_;
  wire _0993_;
  wire _0994_;
  wire _0995_;
  wire _0996_;
  wire _0997_;
  wire _0998_;
  wire _0999_;
  wire _1000_;
  wire _1001_;
  wire _1002_;
  wire _1003_;
  wire _1004_;
  wire _1005_;
  wire _1006_;
  wire _1007_;
  wire _1008_;
  wire _1009_;
  wire _1010_;
  wire _1011_;
  wire _1012_;
  wire _1013_;
  wire _1014_;
  wire _1015_;
  wire _1016_;
  wire _1017_;
  wire _1018_;
  wire _1019_;
  wire _1020_;
  wire _1021_;
  wire _1022_;
  wire _1023_;
  wire _1024_;
  wire _1025_;
  wire _1026_;
  wire _1027_;
  wire _1028_;
  wire _1029_;
  wire _1030_;
  wire _1031_;
  wire _1032_;
  wire _1033_;
  wire _1034_;
  wire _1035_;
  wire _1036_;
  wire _1037_;
  wire _1038_;
  wire _1039_;
  wire _1040_;
  wire _1041_;
  wire _1042_;
  wire _1043_;
  wire _1044_;
  wire _1045_;
  wire _1046_;
  wire _1047_;
  wire _1048_;
  wire _1049_;
  wire _1050_;
  wire _1051_;
  wire _1052_;
  wire _1053_;
  wire _1054_;
  wire _1055_;
  wire _1056_;
  wire _1057_;
  wire _1058_;
  wire _1059_;
  wire _1060_;
  wire _1061_;
  wire _1062_;
  wire _1063_;
  wire _1064_;
  wire _1065_;
  wire _1066_;
  wire _1067_;
  wire _1068_;
  wire _1069_;
  wire _1070_;
  wire _1071_;
  wire _1072_;
  wire _1073_;
  wire _1074_;
  wire _1075_;
  wire _1076_;
  wire _1077_;
  wire _1078_;
  wire _1079_;
  wire _1080_;
  wire _1081_;
  wire _1082_;
  wire _1083_;
  wire _1084_;
  wire _1085_;
  wire _1086_;
  wire _1087_;
  wire _1088_;
  wire _1089_;
  wire _1090_;
  wire _1091_;
  wire _1092_;
  wire _1093_;
  wire _1094_;
  wire _1095_;
  wire _1096_;
  wire _1097_;
  wire _1098_;
  wire _1099_;
  wire _1100_;
  wire _1101_;
  wire _1102_;
  wire _1103_;
  wire _1104_;
  wire _1105_;
  wire _1106_;
  wire _1107_;
  wire _1108_;
  wire _1109_;
  wire _1110_;
  wire _1111_;
  wire _1112_;
  wire _1113_;
  wire _1114_;
  wire _1115_;
  wire _1116_;
  wire _1117_;
  wire _1118_;
  wire _1119_;
  wire _1120_;
  wire _1121_;
  wire _1122_;
  wire _1123_;
  wire _1124_;
  wire _1125_;
  wire _1126_;
  wire _1127_;
  wire _1128_;
  wire _1129_;
  wire _1130_;
  wire _1131_;
  wire _1132_;
  wire _1133_;
  wire _1134_;
  wire _1135_;
  wire _1136_;
  wire _1137_;
  wire _1138_;
  wire _1139_;
  wire _1140_;
  wire _1141_;
  wire _1142_;
  wire _1143_;
  wire _1144_;
  wire _1145_;
  wire _1146_;
  wire _1147_;
  wire _1148_;
  wire _1149_;
  wire _1150_;
  wire _1151_;
  wire _1152_;
  wire _1153_;
  wire _1154_;
  wire _1155_;
  wire _1156_;
  wire _1157_;
  wire _1158_;
  wire _1159_;
  wire _1160_;
  wire _1161_;
  wire _1162_;
  wire _1163_;
  wire _1164_;
  wire _1165_;
  wire _1166_;
  wire _1167_;
  wire _1168_;
  wire _1169_;
  wire _1170_;
  wire _1171_;
  wire _1172_;
  wire _1173_;
  wire _1174_;
  wire _1175_;
  wire _1176_;
  wire _1177_;
  wire _1178_;
  wire _1179_;
  wire _1180_;
  wire _1181_;
  wire _1182_;
  wire _1183_;
  wire _1184_;
  wire _1185_;
  wire _1186_;
  wire _1187_;
  wire _1188_;
  wire _1189_;
  wire _1190_;
  wire _1191_;
  wire _1192_;
  wire _1193_;
  wire _1194_;
  wire _1195_;
  wire _1196_;
  wire _1197_;
  wire _1198_;
  wire _1199_;
  wire _1200_;
  wire _1201_;
  wire _1202_;
  wire _1203_;
  wire _1204_;
  wire _1205_;
  wire _1206_;
  wire _1207_;
  wire _1208_;
  wire _1209_;
  wire _1210_;
  wire _1211_;
  wire _1212_;
  wire _1213_;
  wire _1214_;
  wire _1215_;
  wire _1216_;
  wire _1217_;
  wire _1218_;
  wire _1219_;
  wire _1220_;
  wire _1221_;
  wire _1222_;
  wire _1223_;
  wire _1224_;
  wire _1225_;
  wire _1226_;
  wire _1227_;
  wire _1228_;
  wire _1229_;
  wire _1230_;
  wire _1231_;
  wire _1232_;
  wire _1233_;
  wire _1234_;
  wire _1235_;
  wire _1236_;
  wire _1237_;
  wire _1238_;
  wire _1239_;
  wire _1240_;
  wire _1241_;
  wire _1242_;
  wire _1243_;
  wire _1244_;
  wire _1245_;
  wire _1246_;
  wire _1247_;
  wire _1248_;
  wire _1249_;
  wire _1250_;
  wire _1251_;
  wire _1252_;
  wire _1253_;
  wire _1254_;
  wire _1255_;
  wire _1256_;
  wire _1257_;
  wire _1258_;
  wire _1259_;
  wire _1260_;
  wire _1261_;
  wire _1262_;
  wire _1263_;
  wire _1264_;
  wire _1265_;
  wire _1266_;
  wire _1267_;
  wire _1268_;
  wire _1269_;
  wire _1270_;
  wire _1271_;
  wire _1272_;
  wire _1273_;
  wire _1274_;
  wire _1275_;
  wire _1276_;
  wire _1277_;
  wire _1278_;
  wire _1279_;
  wire _1280_;
  wire _1281_;
  wire _1282_;
  wire _1283_;
  wire _1284_;
  wire _1285_;
  wire _1286_;
  wire _1287_;
  wire _1288_;
  wire _1289_;
  wire _1290_;
  wire _1291_;
  wire _1292_;
  wire _1293_;
  wire _1294_;
  wire _1295_;
  wire _1296_;
  wire _1297_;
  wire _1298_;
  wire _1299_;
  wire _1300_;
  wire _1301_;
  wire _1302_;
  wire _1303_;
  wire _1304_;
  wire _1305_;
  wire _1306_;
  wire _1307_;
  wire _1308_;
  wire _1309_;
  wire _1310_;
  wire _1311_;
  wire _1312_;
  wire _1313_;
  wire _1314_;
  wire _1315_;
  wire _1316_;
  wire _1317_;
  wire _1318_;
  wire _1319_;
  wire _1320_;
  wire _1321_;
  wire _1322_;
  wire _1323_;
  wire _1324_;
  wire _1325_;
  wire _1326_;
  wire _1327_;
  wire _1328_;
  wire _1329_;
  wire _1330_;
  wire _1331_;
  wire _1332_;
  wire _1333_;
  wire _1334_;
  wire _1335_;
  wire _1336_;
  wire _1337_;
  wire _1338_;
  wire _1339_;
  wire _1340_;
  wire _1341_;
  wire _1342_;
  wire _1343_;
  wire _1344_;
  wire _1345_;
  wire _1346_;
  wire _1347_;
  wire _1348_;
  wire _1349_;
  wire _1350_;
  wire _1351_;
  wire _1352_;
  wire _1353_;
  wire _1354_;
  wire _1355_;
  wire _1356_;
  wire _1357_;
  wire _1358_;
  wire _1359_;
  wire _1360_;
  wire _1361_;
  wire _1362_;
  wire _1363_;
  wire _1364_;
  wire _1365_;
  wire _1366_;
  wire _1367_;
  wire _1368_;
  wire _1369_;
  wire _1370_;
  wire _1371_;
  wire _1372_;
  wire _1373_;
  wire _1374_;
  wire _1375_;
  wire _1376_;
  wire _1377_;
  wire _1378_;
  wire _1379_;
  wire _1380_;
  wire _1381_;
  wire _1382_;
  wire _1383_;
  wire _1384_;
  wire _1385_;
  wire _1386_;
  wire _1387_;
  wire _1388_;
  wire _1389_;
  wire _1390_;
  wire _1391_;
  wire _1392_;
  wire _1393_;
  wire _1394_;
  wire _1395_;
  wire _1396_;
  wire _1397_;
  wire _1398_;
  wire _1399_;
  wire _1400_;
  wire _1401_;
  wire _1402_;
  wire _1403_;
  wire _1404_;
  wire _1405_;
  wire _1406_;
  wire _1407_;
  wire _1408_;
  wire _1409_;
  wire _1410_;
  wire _1411_;
  wire _1412_;
  wire _1413_;
  wire _1414_;
  wire _1415_;
  wire _1416_;
  wire _1417_;
  wire _1418_;
  wire _1419_;
  wire _1420_;
  wire _1421_;
  wire _1422_;
  wire _1423_;
  wire _1424_;
  wire _1425_;
  wire _1426_;
  wire _1427_;
  wire _1428_;
  wire _1429_;
  wire _1430_;
  wire _1431_;
  wire _1432_;
  wire _1433_;
  wire _1434_;
  wire _1435_;
  wire _1436_;
  wire _1437_;
  wire _1438_;
  wire _1439_;
  wire _1440_;
  wire _1441_;
  wire _1442_;
  wire _1443_;
  wire _1444_;
  wire _1445_;
  wire _1446_;
  wire _1447_;
  wire _1448_;
  wire _1449_;
  wire _1450_;
  wire _1451_;
  wire _1452_;
  wire _1453_;
  wire _1454_;
  wire _1455_;
  wire _1456_;
  wire _1457_;
  wire _1458_;
  wire _1459_;
  wire _1460_;
  wire _1461_;
  wire _1462_;
  wire _1463_;
  wire _1464_;
  wire _1465_;
  wire _1466_;
  wire _1467_;
  wire _1468_;
  wire _1469_;
  wire _1470_;
  wire _1471_;
  wire _1472_;
  wire _1473_;
  wire _1474_;
  wire _1475_;
  wire _1476_;
  wire _1477_;
  wire _1478_;
  wire _1479_;
  wire _1480_;
  wire _1481_;
  wire _1482_;
  wire _1483_;
  wire _1484_;
  wire _1485_;
  wire _1486_;
  wire _1487_;
  wire _1488_;
  wire _1489_;
  wire _1490_;
  wire _1491_;
  wire _1492_;
  wire _1493_;
  wire _1494_;
  wire _1495_;
  wire _1496_;
  wire _1497_;
  wire _1498_;
  wire _1499_;
  wire _1500_;
  wire _1501_;
  wire _1502_;
  wire _1503_;
  wire _1504_;
  wire _1505_;
  wire _1506_;
  wire _1507_;
  wire _1508_;
  wire _1509_;
  wire _1510_;
  wire _1511_;
  wire _1512_;
  wire _1513_;
  wire _1514_;
  wire _1515_;
  wire _1516_;
  wire _1517_;
  wire _1518_;
  wire _1519_;
  wire _1520_;
  wire _1521_;
  wire _1522_;
  wire _1523_;
  wire _1524_;
  wire _1525_;
  wire _1526_;
  wire _1527_;
  wire _1528_;
  wire _1529_;
  wire _1530_;
  wire _1531_;
  wire _1532_;
  wire _1533_;
  wire _1534_;
  wire _1535_;
  wire _1536_;
  wire _1537_;
  wire _1538_;
  wire _1539_;
  wire _1540_;
  wire _1541_;
  wire _1542_;
  wire _1543_;
  wire _1544_;
  wire _1545_;
  wire _1546_;
  wire _1547_;
  wire _1548_;
  wire _1549_;
  wire _1550_;
  wire _1551_;
  wire _1552_;
  wire _1553_;
  wire _1554_;
  wire _1555_;
  wire _1556_;
  wire _1557_;
  wire _1558_;
  wire _1559_;
  wire _1560_;
  wire _1561_;
  wire _1562_;
  wire _1563_;
  wire _1564_;
  wire _1565_;
  wire _1566_;
  wire _1567_;
  wire _1568_;
  wire _1569_;
  wire _1570_;
  wire _1571_;
  wire _1572_;
  wire _1573_;
  wire _1574_;
  wire _1575_;
  wire _1576_;
  wire _1577_;
  wire _1578_;
  wire _1579_;
  wire _1580_;
  wire _1581_;
  wire _1582_;
  wire _1583_;
  wire _1584_;
  wire _1585_;
  wire _1586_;
  wire _1587_;
  wire _1588_;
  wire _1589_;
  wire _1590_;
  wire _1591_;
  wire _1592_;
  wire _1593_;
  wire _1594_;
  wire _1595_;
  wire _1596_;
  wire _1597_;
  wire _1598_;
  wire _1599_;
  wire [1:0] buffer_head;
  wire [1:0] buffer_tail;
  input clk;
  wire clk;
  input [3:0] dest_addr;
  wire [3:0] dest_addr;
  wire [2:0] network_state;
  wire [63:0] packet_buffer_0;
  wire [63:0] packet_buffer_1;
  wire [63:0] packet_buffer_2;
  wire [63:0] packet_buffer_3;
  wire [3:0] packet_count;
  input [63:0] packet_in;
  wire [63:0] packet_in;
  output [63:0] packet_out;
  wire [63:0] packet_out;
  output packet_ready;
  wire packet_ready;
  input packet_valid;
  wire packet_valid;
  output route_error;
  wire route_error;
  input rst;
  wire rst;
    not _1600_(_0000_, rst);
    not _1601_(_1377_, network_state[2]);
    not _1602_(_1378_, network_state[0]);
    nor _1603_(_1379_, network_state[1], _1378_);
    and _1604_(_1380_, _1379_, _1377_);
    and _1605_(_1381_, _1380_, _0000_);
    and _1606_(_1382_, buffer_tail[1], buffer_tail[0]);
    and _1607_(_1383_, _1382_, _1381_);
    not _1608_(_1384_, _1383_);
    and _1609_(_1385_, _1384_, packet_buffer_3[52]);
    and _1610_(_1386_, _1383_, packet_in[52]);
    or _1611_(_0013_, _1386_, _1385_);
    and _1612_(_1387_, _1384_, packet_buffer_3[53]);
    and _1613_(_1388_, _1383_, packet_in[53]);
    or _1614_(_0014_, _1388_, _1387_);
    and _1615_(_1389_, _1384_, packet_buffer_3[54]);
    and _1616_(_1390_, _1383_, packet_in[54]);
    or _1617_(_0015_, _1390_, _1389_);
    and _1618_(_1391_, _1384_, packet_buffer_3[55]);
    and _1619_(_1392_, _1383_, packet_in[55]);
    or _1620_(_0016_, _1392_, _1391_);
    and _1621_(_1393_, _1384_, packet_buffer_3[56]);
    and _1622_(_1394_, _1383_, packet_in[56]);
    or _1623_(_0017_, _1394_, _1393_);
    and _1624_(_1395_, _1384_, packet_buffer_3[57]);
    and _1625_(_1396_, _1383_, packet_in[57]);
    or _1626_(_0018_, _1396_, _1395_);
    and _1627_(_1397_, _1384_, packet_buffer_3[58]);
    and _1628_(_1398_, _1383_, packet_in[58]);
    or _1629_(_0019_, _1398_, _1397_);
    and _1630_(_1399_, _1384_, packet_buffer_3[59]);
    and _1631_(_1400_, _1383_, packet_in[59]);
    or _1632_(_0020_, _1400_, _1399_);
    and _1633_(_1401_, _1384_, packet_buffer_3[60]);
    and _1634_(_1402_, _1383_, packet_in[60]);
    or _1635_(_0021_, _1402_, _1401_);
    and _1636_(_1403_, _1384_, packet_buffer_3[61]);
    and _1637_(_1404_, _1383_, packet_in[61]);
    or _1638_(_0022_, _1404_, _1403_);
    and _1639_(_1405_, _1384_, packet_buffer_3[62]);
    and _1640_(_1406_, _1383_, packet_in[62]);
    or _1641_(_0023_, _1406_, _1405_);
    and _1642_(_1407_, _1384_, packet_buffer_3[63]);
    and _1643_(_1408_, _1383_, packet_in[63]);
    or _1644_(_0024_, _1408_, _1407_);
    and _1645_(_1409_, network_state[1], network_state[0]);
    and _1646_(_1410_, _1409_, _1377_);
    nor _1647_(_1411_, _1410_, _1380_);
    and _1648_(_1412_, _1411_, packet_count[0]);
    not _1649_(_1413_, _1411_);
    not _1650_(_1414_, packet_count[0]);
    and _1651_(_1415_, _1410_, _1414_);
    and _1652_(_1416_, _1380_, _1414_);
    or _1653_(_1417_, _1416_, _1415_);
    and _1654_(_1418_, _1417_, _1413_);
    or _1655_(_0029_, _1418_, _1412_);
    and _1656_(_1419_, _1411_, packet_count[1]);
    xnor _1657_(_1420_, packet_count[1], packet_count[0]);
    and _1658_(_1421_, _1420_, _1410_);
    xor _1659_(_1422_, packet_count[1], packet_count[0]);
    and _1660_(_1423_, _1422_, _1380_);
    or _1661_(_1424_, _1423_, _1421_);
    and _1662_(_1425_, _1424_, _1413_);
    or _1663_(_0030_, _1425_, _1419_);
    and _1664_(_1426_, _1411_, packet_count[2]);
    nor _1665_(_1427_, packet_count[1], packet_count[0]);
    xor _1666_(_1428_, _1427_, packet_count[2]);
    and _1667_(_1429_, _1428_, _1410_);
    and _1668_(_1430_, packet_count[1], packet_count[0]);
    xor _1669_(_1431_, _1430_, packet_count[2]);
    and _1670_(_1432_, _1431_, _1380_);
    or _1671_(_1433_, _1432_, _1429_);
    and _1672_(_1434_, _1433_, _1413_);
    or _1673_(_0031_, _1434_, _1426_);
    and _1674_(_1435_, _1411_, packet_count[3]);
    not _1675_(_1436_, packet_count[2]);
    and _1676_(_1437_, _1427_, _1436_);
    xor _1677_(_1438_, _1437_, packet_count[3]);
    and _1678_(_1439_, _1438_, _1410_);
    and _1679_(_1440_, _1430_, packet_count[2]);
    xor _1680_(_1441_, _1440_, packet_count[3]);
    and _1681_(_1442_, _1441_, _1380_);
    or _1682_(_1443_, _1442_, _1439_);
    and _1683_(_1444_, _1443_, _1413_);
    or _1684_(_0032_, _1444_, _1435_);
    nor _1685_(_1445_, packet_count[1], packet_count[0]);
    nor _1686_(_1446_, packet_count[3], _1436_);
    nand _1687_(_1447_, _1446_, _1445_);
    and _1688_(_1448_, _1447_, packet_valid);
    nor _1689_(_1449_, network_state[1], network_state[0]);
    and _1690_(_1450_, _1449_, _1377_);
    not _1691_(_1451_, _1450_);
    nor _1692_(_1452_, _1451_, _1448_);
    and _1693_(_1453_, _1452_, network_state[0]);
    not _1694_(_1454_, _1452_);
    nor _1695_(_1455_, packet_count[3], packet_count[2]);
    nand _1696_(_1456_, _1455_, _1445_);
    and _1697_(_1457_, network_state[1], _1378_);
    and _1698_(_1458_, _1457_, _1377_);
    and _1699_(_1459_, _1458_, _1456_);
    and _1700_(_1460_, _1450_, _1448_);
    or _1701_(_1461_, _1460_, _1459_);
    or _1702_(_1462_, _1458_, _1380_);
    or _1703_(_1463_, _1462_, _1450_);
    and _1704_(_1464_, _1463_, _1461_);
    and _1705_(_1465_, _1464_, _1454_);
    or _1706_(_0033_, _1465_, _1453_);
    and _1707_(_1466_, _1452_, network_state[1]);
    or _1708_(_1467_, _1459_, _1380_);
    and _1709_(_1468_, _1467_, _1463_);
    and _1710_(_1469_, _1468_, _1454_);
    or _1711_(_0034_, _1469_, _1466_);
    and _1712_(_0035_, _1452_, network_state[2]);
    and _1713_(_1470_, _1410_, _0000_);
    not _1714_(_1471_, _1470_);
    and _1715_(_1472_, _1471_, packet_out[0]);
    and _1716_(_1473_, buffer_head[1], buffer_head[0]);
    and _1717_(_1474_, _1473_, packet_buffer_3[0]);
    not _1718_(_1475_, buffer_head[1]);
    nor _1719_(_1476_, _1475_, buffer_head[0]);
    and _1720_(_1477_, _1476_, packet_buffer_2[0]);
    or _1721_(_1478_, _1477_, _1474_);
    and _1722_(_1479_, _1475_, buffer_head[0]);
    and _1723_(_1480_, _1479_, packet_buffer_1[0]);
    nor _1724_(_1481_, buffer_head[1], buffer_head[0]);
    and _1725_(_1482_, _1481_, packet_buffer_0[0]);
    or _1726_(_1483_, _1482_, _1480_);
    or _1727_(_1484_, _1483_, _1478_);
    or _1728_(_1485_, _1476_, _1473_);
    or _1729_(_1486_, _1481_, _1479_);
    or _1730_(_1487_, _1486_, _1485_);
    and _1731_(_1488_, _1487_, _1484_);
    and _1732_(_1489_, _1488_, _1470_);
    or _1733_(_0036_, _1489_, _1472_);
    and _1734_(_1490_, _1471_, packet_out[1]);
    and _1735_(_1491_, _1473_, packet_buffer_3[1]);
    and _1736_(_1492_, _1476_, packet_buffer_2[1]);
    or _1737_(_1493_, _1492_, _1491_);
    and _1738_(_1494_, _1479_, packet_buffer_1[1]);
    and _1739_(_1495_, _1481_, packet_buffer_0[1]);
    or _1740_(_1496_, _1495_, _1494_);
    or _1741_(_1497_, _1496_, _1493_);
    and _1742_(_1498_, _1497_, _1487_);
    and _1743_(_1499_, _1498_, _1470_);
    or _1744_(_0037_, _1499_, _1490_);
    and _1745_(_1500_, _1471_, packet_out[2]);
    and _1746_(_1501_, _1473_, packet_buffer_3[2]);
    and _1747_(_1502_, _1476_, packet_buffer_2[2]);
    or _1748_(_1503_, _1502_, _1501_);
    and _1749_(_1504_, _1479_, packet_buffer_1[2]);
    and _1750_(_1505_, _1481_, packet_buffer_0[2]);
    or _1751_(_1506_, _1505_, _1504_);
    or _1752_(_1507_, _1506_, _1503_);
    and _1753_(_1508_, _1507_, _1487_);
    and _1754_(_1509_, _1508_, _1470_);
    or _1755_(_0038_, _1509_, _1500_);
    and _1756_(_1510_, _1471_, packet_out[3]);
    and _1757_(_1511_, _1473_, packet_buffer_3[3]);
    and _1758_(_1512_, _1476_, packet_buffer_2[3]);
    or _1759_(_1513_, _1512_, _1511_);
    and _1760_(_1514_, _1479_, packet_buffer_1[3]);
    and _1761_(_1515_, _1481_, packet_buffer_0[3]);
    or _1762_(_1516_, _1515_, _1514_);
    or _1763_(_1517_, _1516_, _1513_);
    and _1764_(_1518_, _1517_, _1487_);
    and _1765_(_1519_, _1518_, _1470_);
    or _1766_(_0039_, _1519_, _1510_);
    and _1767_(_1520_, _1471_, packet_out[4]);
    and _1768_(_1521_, _1473_, packet_buffer_3[4]);
    and _1769_(_1522_, _1476_, packet_buffer_2[4]);
    or _1770_(_1523_, _1522_, _1521_);
    and _1771_(_1524_, _1479_, packet_buffer_1[4]);
    and _1772_(_1525_, _1481_, packet_buffer_0[4]);
    or _1773_(_1526_, _1525_, _1524_);
    or _1774_(_1527_, _1526_, _1523_);
    and _1775_(_1528_, _1527_, _1487_);
    and _1776_(_1529_, _1528_, _1470_);
    or _1777_(_0040_, _1529_, _1520_);
    and _1778_(_1530_, _1471_, packet_out[5]);
    and _1779_(_1531_, _1473_, packet_buffer_3[5]);
    and _1780_(_1532_, _1476_, packet_buffer_2[5]);
    or _1781_(_1533_, _1532_, _1531_);
    and _1782_(_1534_, _1479_, packet_buffer_1[5]);
    and _1783_(_1535_, _1481_, packet_buffer_0[5]);
    or _1784_(_1536_, _1535_, _1534_);
    or _1785_(_1537_, _1536_, _1533_);
    and _1786_(_1538_, _1537_, _1487_);
    and _1787_(_1539_, _1538_, _1470_);
    or _1788_(_0041_, _1539_, _1530_);
    and _1789_(_1540_, _1471_, packet_out[6]);
    and _1790_(_1541_, _1473_, packet_buffer_3[6]);
    and _1791_(_1542_, _1476_, packet_buffer_2[6]);
    or _1792_(_1543_, _1542_, _1541_);
    and _1793_(_1544_, _1479_, packet_buffer_1[6]);
    and _1794_(_1545_, _1481_, packet_buffer_0[6]);
    or _1795_(_1546_, _1545_, _1544_);
    or _1796_(_1547_, _1546_, _1543_);
    and _1797_(_1548_, _1547_, _1487_);
    and _1798_(_1549_, _1548_, _1470_);
    or _1799_(_0042_, _1549_, _1540_);
    and _1800_(_1550_, _1471_, packet_out[7]);
    and _1801_(_1551_, _1473_, packet_buffer_3[7]);
    and _1802_(_1552_, _1476_, packet_buffer_2[7]);
    or _1803_(_1553_, _1552_, _1551_);
    and _1804_(_1554_, _1479_, packet_buffer_1[7]);
    and _1805_(_1555_, _1481_, packet_buffer_0[7]);
    or _1806_(_1556_, _1555_, _1554_);
    or _1807_(_1557_, _1556_, _1553_);
    and _1808_(_1558_, _1557_, _1487_);
    and _1809_(_1559_, _1558_, _1470_);
    or _1810_(_0043_, _1559_, _1550_);
    and _1811_(_1560_, _1471_, packet_out[8]);
    and _1812_(_1561_, _1473_, packet_buffer_3[8]);
    and _1813_(_1562_, _1476_, packet_buffer_2[8]);
    or _1814_(_1563_, _1562_, _1561_);
    and _1815_(_1564_, _1479_, packet_buffer_1[8]);
    and _1816_(_1565_, _1481_, packet_buffer_0[8]);
    or _1817_(_1566_, _1565_, _1564_);
    or _1818_(_1567_, _1566_, _1563_);
    and _1819_(_1568_, _1567_, _1487_);
    and _1820_(_1569_, _1568_, _1470_);
    or _1821_(_0044_, _1569_, _1560_);
    and _1822_(_1570_, _1471_, packet_out[9]);
    and _1823_(_1571_, _1473_, packet_buffer_3[9]);
    and _1824_(_1572_, _1476_, packet_buffer_2[9]);
    or _1825_(_1573_, _1572_, _1571_);
    and _1826_(_1574_, _1479_, packet_buffer_1[9]);
    and _1827_(_1575_, _1481_, packet_buffer_0[9]);
    or _1828_(_1576_, _1575_, _1574_);
    or _1829_(_1577_, _1576_, _1573_);
    and _1830_(_1578_, _1577_, _1487_);
    and _1831_(_1579_, _1578_, _1470_);
    or _1832_(_0045_, _1579_, _1570_);
    and _1833_(_1580_, _1471_, packet_out[10]);
    and _1834_(_1581_, _1473_, packet_buffer_3[10]);
    and _1835_(_1582_, _1476_, packet_buffer_2[10]);
    or _1836_(_1583_, _1582_, _1581_);
    and _1837_(_1584_, _1479_, packet_buffer_1[10]);
    and _1838_(_1585_, _1481_, packet_buffer_0[10]);
    or _1839_(_1586_, _1585_, _1584_);
    or _1840_(_1587_, _1586_, _1583_);
    and _1841_(_1588_, _1587_, _1487_);
    and _1842_(_1589_, _1588_, _1470_);
    or _1843_(_0046_, _1589_, _1580_);
    and _1844_(_1590_, _1471_, packet_out[11]);
    and _1845_(_1591_, _1473_, packet_buffer_3[11]);
    and _1846_(_1592_, _1476_, packet_buffer_2[11]);
    or _1847_(_1593_, _1592_, _1591_);
    and _1848_(_1594_, _1479_, packet_buffer_1[11]);
    and _1849_(_1595_, _1481_, packet_buffer_0[11]);
    or _1850_(_1596_, _1595_, _1594_);
    or _1851_(_1597_, _1596_, _1593_);
    and _1852_(_1598_, _1597_, _1487_);
    and _1853_(_1599_, _1598_, _1470_);
    or _1854_(_0047_, _1599_, _1590_);
    and _1855_(_0346_, _1471_, packet_out[12]);
    and _1856_(_0347_, _1473_, packet_buffer_3[12]);
    and _1857_(_0348_, _1476_, packet_buffer_2[12]);
    or _1858_(_0349_, _0348_, _0347_);
    and _1859_(_0350_, _1479_, packet_buffer_1[12]);
    and _1860_(_0351_, _1481_, packet_buffer_0[12]);
    or _1861_(_0352_, _0351_, _0350_);
    or _1862_(_0353_, _0352_, _0349_);
    and _1863_(_0354_, _0353_, _1487_);
    and _1864_(_0355_, _0354_, _1470_);
    or _1865_(_0048_, _0355_, _0346_);
    and _1866_(_0356_, _1471_, packet_out[13]);
    and _1867_(_0357_, _1473_, packet_buffer_3[13]);
    and _1868_(_0358_, _1476_, packet_buffer_2[13]);
    or _1869_(_0359_, _0358_, _0357_);
    and _1870_(_0360_, _1479_, packet_buffer_1[13]);
    and _1871_(_0361_, _1481_, packet_buffer_0[13]);
    or _1872_(_0362_, _0361_, _0360_);
    or _1873_(_0363_, _0362_, _0359_);
    and _1874_(_0364_, _0363_, _1487_);
    and _1875_(_0365_, _0364_, _1470_);
    or _1876_(_0049_, _0365_, _0356_);
    and _1877_(_0366_, _1471_, packet_out[14]);
    and _1878_(_0367_, _1473_, packet_buffer_3[14]);
    and _1879_(_0368_, _1476_, packet_buffer_2[14]);
    or _1880_(_0369_, _0368_, _0367_);
    and _1881_(_0370_, _1479_, packet_buffer_1[14]);
    and _1882_(_0371_, _1481_, packet_buffer_0[14]);
    or _1883_(_0372_, _0371_, _0370_);
    or _1884_(_0373_, _0372_, _0369_);
    and _1885_(_0374_, _0373_, _1487_);
    and _1886_(_0375_, _0374_, _1470_);
    or _1887_(_0050_, _0375_, _0366_);
    and _1888_(_0376_, _1471_, packet_out[15]);
    and _1889_(_0377_, _1473_, packet_buffer_3[15]);
    and _1890_(_0378_, _1476_, packet_buffer_2[15]);
    or _1891_(_0379_, _0378_, _0377_);
    and _1892_(_0380_, _1479_, packet_buffer_1[15]);
    and _1893_(_0381_, _1481_, packet_buffer_0[15]);
    or _1894_(_0382_, _0381_, _0380_);
    or _1895_(_0383_, _0382_, _0379_);
    and _1896_(_0384_, _0383_, _1487_);
    and _1897_(_0385_, _0384_, _1470_);
    or _1898_(_0051_, _0385_, _0376_);
    and _1899_(_0386_, _1471_, packet_out[16]);
    and _1900_(_0387_, _1473_, packet_buffer_3[16]);
    and _1901_(_0388_, _1476_, packet_buffer_2[16]);
    or _1902_(_0389_, _0388_, _0387_);
    and _1903_(_0390_, _1479_, packet_buffer_1[16]);
    and _1904_(_0391_, _1481_, packet_buffer_0[16]);
    or _1905_(_0392_, _0391_, _0390_);
    or _1906_(_0393_, _0392_, _0389_);
    and _1907_(_0394_, _0393_, _1487_);
    and _1908_(_0395_, _0394_, _1470_);
    or _1909_(_0052_, _0395_, _0386_);
    and _1910_(_0396_, _1471_, packet_out[17]);
    and _1911_(_0397_, _1473_, packet_buffer_3[17]);
    and _1912_(_0398_, _1476_, packet_buffer_2[17]);
    or _1913_(_0399_, _0398_, _0397_);
    and _1914_(_0400_, _1479_, packet_buffer_1[17]);
    and _1915_(_0401_, _1481_, packet_buffer_0[17]);
    or _1916_(_0402_, _0401_, _0400_);
    or _1917_(_0403_, _0402_, _0399_);
    and _1918_(_0404_, _0403_, _1487_);
    and _1919_(_0405_, _0404_, _1470_);
    or _1920_(_0053_, _0405_, _0396_);
    and _1921_(_0406_, _1471_, packet_out[18]);
    and _1922_(_0407_, _1473_, packet_buffer_3[18]);
    and _1923_(_0408_, _1476_, packet_buffer_2[18]);
    or _1924_(_0409_, _0408_, _0407_);
    and _1925_(_0410_, _1479_, packet_buffer_1[18]);
    and _1926_(_0411_, _1481_, packet_buffer_0[18]);
    or _1927_(_0412_, _0411_, _0410_);
    or _1928_(_0413_, _0412_, _0409_);
    and _1929_(_0414_, _0413_, _1487_);
    and _1930_(_0415_, _0414_, _1470_);
    or _1931_(_0054_, _0415_, _0406_);
    and _1932_(_0416_, _1471_, packet_out[19]);
    and _1933_(_0417_, _1473_, packet_buffer_3[19]);
    and _1934_(_0418_, _1476_, packet_buffer_2[19]);
    or _1935_(_0419_, _0418_, _0417_);
    and _1936_(_0420_, _1479_, packet_buffer_1[19]);
    and _1937_(_0421_, _1481_, packet_buffer_0[19]);
    or _1938_(_0422_, _0421_, _0420_);
    or _1939_(_0423_, _0422_, _0419_);
    and _1940_(_0424_, _0423_, _1487_);
    and _1941_(_0425_, _0424_, _1470_);
    or _1942_(_0055_, _0425_, _0416_);
    and _1943_(_0426_, _1471_, packet_out[20]);
    and _1944_(_0427_, _1473_, packet_buffer_3[20]);
    and _1945_(_0428_, _1476_, packet_buffer_2[20]);
    or _1946_(_0429_, _0428_, _0427_);
    and _1947_(_0430_, _1479_, packet_buffer_1[20]);
    and _1948_(_0431_, _1481_, packet_buffer_0[20]);
    or _1949_(_0432_, _0431_, _0430_);
    or _1950_(_0433_, _0432_, _0429_);
    and _1951_(_0434_, _0433_, _1487_);
    and _1952_(_0435_, _0434_, _1470_);
    or _1953_(_0056_, _0435_, _0426_);
    and _1954_(_0436_, _1471_, packet_out[21]);
    and _1955_(_0437_, _1473_, packet_buffer_3[21]);
    and _1956_(_0438_, _1476_, packet_buffer_2[21]);
    or _1957_(_0439_, _0438_, _0437_);
    and _1958_(_0440_, _1479_, packet_buffer_1[21]);
    and _1959_(_0441_, _1481_, packet_buffer_0[21]);
    or _1960_(_0442_, _0441_, _0440_);
    or _1961_(_0443_, _0442_, _0439_);
    and _1962_(_0444_, _0443_, _1487_);
    and _1963_(_0445_, _0444_, _1470_);
    or _1964_(_0057_, _0445_, _0436_);
    and _1965_(_0446_, _1471_, packet_out[22]);
    and _1966_(_0447_, _1473_, packet_buffer_3[22]);
    and _1967_(_0448_, _1476_, packet_buffer_2[22]);
    or _1968_(_0449_, _0448_, _0447_);
    and _1969_(_0450_, _1479_, packet_buffer_1[22]);
    and _1970_(_0451_, _1481_, packet_buffer_0[22]);
    or _1971_(_0452_, _0451_, _0450_);
    or _1972_(_0453_, _0452_, _0449_);
    and _1973_(_0454_, _0453_, _1487_);
    and _1974_(_0455_, _0454_, _1470_);
    or _1975_(_0058_, _0455_, _0446_);
    and _1976_(_0456_, _1471_, packet_out[23]);
    and _1977_(_0457_, _1473_, packet_buffer_3[23]);
    and _1978_(_0458_, _1476_, packet_buffer_2[23]);
    or _1979_(_0459_, _0458_, _0457_);
    and _1980_(_0460_, _1479_, packet_buffer_1[23]);
    and _1981_(_0461_, _1481_, packet_buffer_0[23]);
    or _1982_(_0462_, _0461_, _0460_);
    or _1983_(_0463_, _0462_, _0459_);
    and _1984_(_0464_, _0463_, _1487_);
    and _1985_(_0465_, _0464_, _1470_);
    or _1986_(_0059_, _0465_, _0456_);
    and _1987_(_0466_, _1471_, packet_out[24]);
    and _1988_(_0467_, _1473_, packet_buffer_3[24]);
    and _1989_(_0468_, _1476_, packet_buffer_2[24]);
    or _1990_(_0469_, _0468_, _0467_);
    and _1991_(_0470_, _1479_, packet_buffer_1[24]);
    and _1992_(_0471_, _1481_, packet_buffer_0[24]);
    or _1993_(_0472_, _0471_, _0470_);
    or _1994_(_0473_, _0472_, _0469_);
    and _1995_(_0474_, _0473_, _1487_);
    and _1996_(_0475_, _0474_, _1470_);
    or _1997_(_0060_, _0475_, _0466_);
    and _1998_(_0476_, _1471_, packet_out[25]);
    and _1999_(_0477_, _1473_, packet_buffer_3[25]);
    and _2000_(_0478_, _1476_, packet_buffer_2[25]);
    or _2001_(_0479_, _0478_, _0477_);
    and _2002_(_0480_, _1479_, packet_buffer_1[25]);
    and _2003_(_0481_, _1481_, packet_buffer_0[25]);
    or _2004_(_0482_, _0481_, _0480_);
    or _2005_(_0483_, _0482_, _0479_);
    and _2006_(_0484_, _0483_, _1487_);
    and _2007_(_0485_, _0484_, _1470_);
    or _2008_(_0061_, _0485_, _0476_);
    and _2009_(_0486_, _1471_, packet_out[26]);
    and _2010_(_0487_, _1473_, packet_buffer_3[26]);
    and _2011_(_0488_, _1476_, packet_buffer_2[26]);
    or _2012_(_0489_, _0488_, _0487_);
    and _2013_(_0490_, _1479_, packet_buffer_1[26]);
    and _2014_(_0491_, _1481_, packet_buffer_0[26]);
    or _2015_(_0492_, _0491_, _0490_);
    or _2016_(_0493_, _0492_, _0489_);
    and _2017_(_0494_, _0493_, _1487_);
    and _2018_(_0495_, _0494_, _1470_);
    or _2019_(_0062_, _0495_, _0486_);
    and _2020_(_0496_, _1471_, packet_out[27]);
    and _2021_(_0497_, _1473_, packet_buffer_3[27]);
    and _2022_(_0498_, _1476_, packet_buffer_2[27]);
    or _2023_(_0499_, _0498_, _0497_);
    and _2024_(_0500_, _1479_, packet_buffer_1[27]);
    and _2025_(_0501_, _1481_, packet_buffer_0[27]);
    or _2026_(_0502_, _0501_, _0500_);
    or _2027_(_0503_, _0502_, _0499_);
    and _2028_(_0504_, _0503_, _1487_);
    and _2029_(_0505_, _0504_, _1470_);
    or _2030_(_0063_, _0505_, _0496_);
    and _2031_(_0506_, _1471_, packet_out[28]);
    and _2032_(_0507_, _1473_, packet_buffer_3[28]);
    and _2033_(_0508_, _1476_, packet_buffer_2[28]);
    or _2034_(_0509_, _0508_, _0507_);
    and _2035_(_0510_, _1479_, packet_buffer_1[28]);
    and _2036_(_0511_, _1481_, packet_buffer_0[28]);
    or _2037_(_0512_, _0511_, _0510_);
    or _2038_(_0513_, _0512_, _0509_);
    and _2039_(_0514_, _0513_, _1487_);
    and _2040_(_0515_, _0514_, _1470_);
    or _2041_(_0064_, _0515_, _0506_);
    and _2042_(_0516_, _1471_, packet_out[29]);
    and _2043_(_0517_, _1473_, packet_buffer_3[29]);
    and _2044_(_0518_, _1476_, packet_buffer_2[29]);
    or _2045_(_0519_, _0518_, _0517_);
    and _2046_(_0520_, _1479_, packet_buffer_1[29]);
    and _2047_(_0521_, _1481_, packet_buffer_0[29]);
    or _2048_(_0522_, _0521_, _0520_);
    or _2049_(_0523_, _0522_, _0519_);
    and _2050_(_0524_, _0523_, _1487_);
    and _2051_(_0525_, _0524_, _1470_);
    or _2052_(_0065_, _0525_, _0516_);
    and _2053_(_0526_, _1471_, packet_out[30]);
    and _2054_(_0527_, _1473_, packet_buffer_3[30]);
    and _2055_(_0528_, _1476_, packet_buffer_2[30]);
    or _2056_(_0529_, _0528_, _0527_);
    and _2057_(_0530_, _1479_, packet_buffer_1[30]);
    and _2058_(_0531_, _1481_, packet_buffer_0[30]);
    or _2059_(_0532_, _0531_, _0530_);
    or _2060_(_0533_, _0532_, _0529_);
    and _2061_(_0534_, _0533_, _1487_);
    and _2062_(_0535_, _0534_, _1470_);
    or _2063_(_0066_, _0535_, _0526_);
    and _2064_(_0536_, _1471_, packet_out[31]);
    and _2065_(_0537_, _1473_, packet_buffer_3[31]);
    and _2066_(_0538_, _1476_, packet_buffer_2[31]);
    or _2067_(_0539_, _0538_, _0537_);
    and _2068_(_0540_, _1479_, packet_buffer_1[31]);
    and _2069_(_0541_, _1481_, packet_buffer_0[31]);
    or _2070_(_0542_, _0541_, _0540_);
    or _2071_(_0543_, _0542_, _0539_);
    and _2072_(_0544_, _0543_, _1487_);
    and _2073_(_0545_, _0544_, _1470_);
    or _2074_(_0067_, _0545_, _0536_);
    and _2075_(_0546_, _1471_, packet_out[32]);
    and _2076_(_0547_, _1473_, packet_buffer_3[32]);
    and _2077_(_0548_, _1476_, packet_buffer_2[32]);
    or _2078_(_0549_, _0548_, _0547_);
    and _2079_(_0550_, _1479_, packet_buffer_1[32]);
    and _2080_(_0551_, _1481_, packet_buffer_0[32]);
    or _2081_(_0552_, _0551_, _0550_);
    or _2082_(_0553_, _0552_, _0549_);
    and _2083_(_0554_, _0553_, _1487_);
    and _2084_(_0555_, _0554_, _1470_);
    or _2085_(_0068_, _0555_, _0546_);
    and _2086_(_0556_, _1471_, packet_out[33]);
    and _2087_(_0557_, _1473_, packet_buffer_3[33]);
    and _2088_(_0558_, _1476_, packet_buffer_2[33]);
    or _2089_(_0559_, _0558_, _0557_);
    and _2090_(_0560_, _1479_, packet_buffer_1[33]);
    and _2091_(_0561_, _1481_, packet_buffer_0[33]);
    or _2092_(_0562_, _0561_, _0560_);
    or _2093_(_0563_, _0562_, _0559_);
    and _2094_(_0564_, _0563_, _1487_);
    and _2095_(_0565_, _0564_, _1470_);
    or _2096_(_0069_, _0565_, _0556_);
    and _2097_(_0566_, _1471_, packet_out[34]);
    and _2098_(_0567_, _1473_, packet_buffer_3[34]);
    and _2099_(_0568_, _1476_, packet_buffer_2[34]);
    or _2100_(_0569_, _0568_, _0567_);
    and _2101_(_0570_, _1479_, packet_buffer_1[34]);
    and _2102_(_0571_, _1481_, packet_buffer_0[34]);
    or _2103_(_0572_, _0571_, _0570_);
    or _2104_(_0573_, _0572_, _0569_);
    and _2105_(_0574_, _0573_, _1487_);
    and _2106_(_0575_, _0574_, _1470_);
    or _2107_(_0070_, _0575_, _0566_);
    and _2108_(_0576_, _1471_, packet_out[35]);
    and _2109_(_0577_, _1473_, packet_buffer_3[35]);
    and _2110_(_0578_, _1476_, packet_buffer_2[35]);
    or _2111_(_0579_, _0578_, _0577_);
    and _2112_(_0580_, _1479_, packet_buffer_1[35]);
    and _2113_(_0581_, _1481_, packet_buffer_0[35]);
    or _2114_(_0582_, _0581_, _0580_);
    or _2115_(_0583_, _0582_, _0579_);
    and _2116_(_0584_, _0583_, _1487_);
    and _2117_(_0585_, _0584_, _1470_);
    or _2118_(_0071_, _0585_, _0576_);
    and _2119_(_0586_, _1471_, packet_out[36]);
    and _2120_(_0587_, _1473_, packet_buffer_3[36]);
    and _2121_(_0588_, _1476_, packet_buffer_2[36]);
    or _2122_(_0589_, _0588_, _0587_);
    and _2123_(_0590_, _1479_, packet_buffer_1[36]);
    and _2124_(_0591_, _1481_, packet_buffer_0[36]);
    or _2125_(_0592_, _0591_, _0590_);
    or _2126_(_0593_, _0592_, _0589_);
    and _2127_(_0594_, _0593_, _1487_);
    and _2128_(_0595_, _0594_, _1470_);
    or _2129_(_0072_, _0595_, _0586_);
    and _2130_(_0596_, _1471_, packet_out[37]);
    and _2131_(_0597_, _1473_, packet_buffer_3[37]);
    and _2132_(_0598_, _1476_, packet_buffer_2[37]);
    or _2133_(_0599_, _0598_, _0597_);
    and _2134_(_0600_, _1479_, packet_buffer_1[37]);
    and _2135_(_0601_, _1481_, packet_buffer_0[37]);
    or _2136_(_0602_, _0601_, _0600_);
    or _2137_(_0603_, _0602_, _0599_);
    and _2138_(_0604_, _0603_, _1487_);
    and _2139_(_0605_, _0604_, _1470_);
    or _2140_(_0073_, _0605_, _0596_);
    and _2141_(_0606_, _1471_, packet_out[38]);
    and _2142_(_0607_, _1473_, packet_buffer_3[38]);
    and _2143_(_0608_, _1476_, packet_buffer_2[38]);
    or _2144_(_0609_, _0608_, _0607_);
    and _2145_(_0610_, _1479_, packet_buffer_1[38]);
    and _2146_(_0611_, _1481_, packet_buffer_0[38]);
    or _2147_(_0612_, _0611_, _0610_);
    or _2148_(_0613_, _0612_, _0609_);
    and _2149_(_0614_, _0613_, _1487_);
    and _2150_(_0615_, _0614_, _1470_);
    or _2151_(_0074_, _0615_, _0606_);
    and _2152_(_0616_, _1471_, packet_out[39]);
    and _2153_(_0617_, _1473_, packet_buffer_3[39]);
    and _2154_(_0618_, _1476_, packet_buffer_2[39]);
    or _2155_(_0619_, _0618_, _0617_);
    and _2156_(_0620_, _1479_, packet_buffer_1[39]);
    and _2157_(_0621_, _1481_, packet_buffer_0[39]);
    or _2158_(_0622_, _0621_, _0620_);
    or _2159_(_0623_, _0622_, _0619_);
    and _2160_(_0624_, _0623_, _1487_);
    and _2161_(_0625_, _0624_, _1470_);
    or _2162_(_0075_, _0625_, _0616_);
    and _2163_(_0626_, _1471_, packet_out[40]);
    and _2164_(_0627_, _1473_, packet_buffer_3[40]);
    and _2165_(_0628_, _1476_, packet_buffer_2[40]);
    or _2166_(_0629_, _0628_, _0627_);
    and _2167_(_0630_, _1479_, packet_buffer_1[40]);
    and _2168_(_0631_, _1481_, packet_buffer_0[40]);
    or _2169_(_0632_, _0631_, _0630_);
    or _2170_(_0633_, _0632_, _0629_);
    and _2171_(_0634_, _0633_, _1487_);
    and _2172_(_0635_, _0634_, _1470_);
    or _2173_(_0076_, _0635_, _0626_);
    and _2174_(_0636_, _1471_, packet_out[41]);
    and _2175_(_0637_, _1473_, packet_buffer_3[41]);
    and _2176_(_0638_, _1476_, packet_buffer_2[41]);
    or _2177_(_0639_, _0638_, _0637_);
    and _2178_(_0640_, _1479_, packet_buffer_1[41]);
    and _2179_(_0641_, _1481_, packet_buffer_0[41]);
    or _2180_(_0642_, _0641_, _0640_);
    or _2181_(_0643_, _0642_, _0639_);
    and _2182_(_0644_, _0643_, _1487_);
    and _2183_(_0645_, _0644_, _1470_);
    or _2184_(_0077_, _0645_, _0636_);
    and _2185_(_0646_, _1471_, packet_out[42]);
    and _2186_(_0647_, _1473_, packet_buffer_3[42]);
    and _2187_(_0648_, _1476_, packet_buffer_2[42]);
    or _2188_(_0649_, _0648_, _0647_);
    and _2189_(_0650_, _1479_, packet_buffer_1[42]);
    and _2190_(_0651_, _1481_, packet_buffer_0[42]);
    or _2191_(_0652_, _0651_, _0650_);
    or _2192_(_0653_, _0652_, _0649_);
    and _2193_(_0654_, _0653_, _1487_);
    and _2194_(_0655_, _0654_, _1470_);
    or _2195_(_0078_, _0655_, _0646_);
    and _2196_(_0656_, _1471_, packet_out[43]);
    and _2197_(_0657_, _1473_, packet_buffer_3[43]);
    and _2198_(_0658_, _1476_, packet_buffer_2[43]);
    or _2199_(_0659_, _0658_, _0657_);
    and _2200_(_0660_, _1479_, packet_buffer_1[43]);
    and _2201_(_0661_, _1481_, packet_buffer_0[43]);
    or _2202_(_0662_, _0661_, _0660_);
    or _2203_(_0663_, _0662_, _0659_);
    and _2204_(_0664_, _0663_, _1487_);
    and _2205_(_0665_, _0664_, _1470_);
    or _2206_(_0079_, _0665_, _0656_);
    and _2207_(_0666_, _1471_, packet_out[44]);
    and _2208_(_0667_, _1473_, packet_buffer_3[44]);
    and _2209_(_0668_, _1476_, packet_buffer_2[44]);
    or _2210_(_0669_, _0668_, _0667_);
    and _2211_(_0670_, _1479_, packet_buffer_1[44]);
    and _2212_(_0671_, _1481_, packet_buffer_0[44]);
    or _2213_(_0672_, _0671_, _0670_);
    or _2214_(_0673_, _0672_, _0669_);
    and _2215_(_0674_, _0673_, _1487_);
    and _2216_(_0675_, _0674_, _1470_);
    or _2217_(_0080_, _0675_, _0666_);
    and _2218_(_0676_, _1471_, packet_out[45]);
    and _2219_(_0677_, _1473_, packet_buffer_3[45]);
    and _2220_(_0678_, _1476_, packet_buffer_2[45]);
    or _2221_(_0679_, _0678_, _0677_);
    and _2222_(_0680_, _1479_, packet_buffer_1[45]);
    and _2223_(_0681_, _1481_, packet_buffer_0[45]);
    or _2224_(_0682_, _0681_, _0680_);
    or _2225_(_0683_, _0682_, _0679_);
    and _2226_(_0684_, _0683_, _1487_);
    and _2227_(_0685_, _0684_, _1470_);
    or _2228_(_0081_, _0685_, _0676_);
    and _2229_(_0686_, _1471_, packet_out[46]);
    and _2230_(_0687_, _1473_, packet_buffer_3[46]);
    and _2231_(_0688_, _1476_, packet_buffer_2[46]);
    or _2232_(_0689_, _0688_, _0687_);
    and _2233_(_0690_, _1479_, packet_buffer_1[46]);
    and _2234_(_0691_, _1481_, packet_buffer_0[46]);
    or _2235_(_0692_, _0691_, _0690_);
    or _2236_(_0693_, _0692_, _0689_);
    and _2237_(_0694_, _0693_, _1487_);
    and _2238_(_0695_, _0694_, _1470_);
    or _2239_(_0082_, _0695_, _0686_);
    and _2240_(_0696_, _1471_, packet_out[47]);
    and _2241_(_0697_, _1473_, packet_buffer_3[47]);
    and _2242_(_0698_, _1476_, packet_buffer_2[47]);
    or _2243_(_0699_, _0698_, _0697_);
    and _2244_(_0700_, _1479_, packet_buffer_1[47]);
    and _2245_(_0701_, _1481_, packet_buffer_0[47]);
    or _2246_(_0702_, _0701_, _0700_);
    or _2247_(_0703_, _0702_, _0699_);
    and _2248_(_0704_, _0703_, _1487_);
    and _2249_(_0705_, _0704_, _1470_);
    or _2250_(_0083_, _0705_, _0696_);
    and _2251_(_0706_, _1471_, packet_out[48]);
    and _2252_(_0707_, _1473_, packet_buffer_3[48]);
    and _2253_(_0708_, _1476_, packet_buffer_2[48]);
    or _2254_(_0709_, _0708_, _0707_);
    and _2255_(_0710_, _1479_, packet_buffer_1[48]);
    and _2256_(_0711_, _1481_, packet_buffer_0[48]);
    or _2257_(_0712_, _0711_, _0710_);
    or _2258_(_0713_, _0712_, _0709_);
    and _2259_(_0714_, _0713_, _1487_);
    and _2260_(_0715_, _0714_, _1470_);
    or _2261_(_0084_, _0715_, _0706_);
    and _2262_(_0716_, _1471_, packet_out[49]);
    and _2263_(_0717_, _1473_, packet_buffer_3[49]);
    and _2264_(_0718_, _1476_, packet_buffer_2[49]);
    or _2265_(_0719_, _0718_, _0717_);
    and _2266_(_0720_, _1479_, packet_buffer_1[49]);
    and _2267_(_0721_, _1481_, packet_buffer_0[49]);
    or _2268_(_0722_, _0721_, _0720_);
    or _2269_(_0723_, _0722_, _0719_);
    and _2270_(_0724_, _0723_, _1487_);
    and _2271_(_0725_, _0724_, _1470_);
    or _2272_(_0085_, _0725_, _0716_);
    and _2273_(_0726_, _1471_, packet_out[50]);
    and _2274_(_0727_, _1473_, packet_buffer_3[50]);
    and _2275_(_0728_, _1476_, packet_buffer_2[50]);
    or _2276_(_0729_, _0728_, _0727_);
    and _2277_(_0730_, _1479_, packet_buffer_1[50]);
    and _2278_(_0731_, _1481_, packet_buffer_0[50]);
    or _2279_(_0732_, _0731_, _0730_);
    or _2280_(_0733_, _0732_, _0729_);
    and _2281_(_0734_, _0733_, _1487_);
    and _2282_(_0735_, _0734_, _1470_);
    or _2283_(_0086_, _0735_, _0726_);
    and _2284_(_0736_, _1471_, packet_out[51]);
    and _2285_(_0737_, _1473_, packet_buffer_3[51]);
    and _2286_(_0738_, _1476_, packet_buffer_2[51]);
    or _2287_(_0739_, _0738_, _0737_);
    and _2288_(_0740_, _1479_, packet_buffer_1[51]);
    and _2289_(_0741_, _1481_, packet_buffer_0[51]);
    or _2290_(_0742_, _0741_, _0740_);
    or _2291_(_0743_, _0742_, _0739_);
    and _2292_(_0744_, _0743_, _1487_);
    and _2293_(_0745_, _0744_, _1470_);
    or _2294_(_0087_, _0745_, _0736_);
    and _2295_(_0746_, _1471_, packet_out[52]);
    and _2296_(_0747_, _1473_, packet_buffer_3[52]);
    and _2297_(_0748_, _1476_, packet_buffer_2[52]);
    or _2298_(_0749_, _0748_, _0747_);
    and _2299_(_0750_, _1479_, packet_buffer_1[52]);
    and _2300_(_0751_, _1481_, packet_buffer_0[52]);
    or _2301_(_0752_, _0751_, _0750_);
    or _2302_(_0753_, _0752_, _0749_);
    and _2303_(_0754_, _0753_, _1487_);
    and _2304_(_0755_, _0754_, _1470_);
    or _2305_(_0088_, _0755_, _0746_);
    and _2306_(_0756_, _1471_, packet_out[53]);
    and _2307_(_0757_, _1473_, packet_buffer_3[53]);
    and _2308_(_0758_, _1476_, packet_buffer_2[53]);
    or _2309_(_0759_, _0758_, _0757_);
    and _2310_(_0760_, _1479_, packet_buffer_1[53]);
    and _2311_(_0761_, _1481_, packet_buffer_0[53]);
    or _2312_(_0762_, _0761_, _0760_);
    or _2313_(_0763_, _0762_, _0759_);
    and _2314_(_0764_, _0763_, _1487_);
    and _2315_(_0765_, _0764_, _1470_);
    or _2316_(_0089_, _0765_, _0756_);
    and _2317_(_0766_, _1471_, packet_out[54]);
    and _2318_(_0767_, _1473_, packet_buffer_3[54]);
    and _2319_(_0768_, _1476_, packet_buffer_2[54]);
    or _2320_(_0769_, _0768_, _0767_);
    and _2321_(_0770_, _1479_, packet_buffer_1[54]);
    and _2322_(_0771_, _1481_, packet_buffer_0[54]);
    or _2323_(_0772_, _0771_, _0770_);
    or _2324_(_0773_, _0772_, _0769_);
    and _2325_(_0774_, _0773_, _1487_);
    and _2326_(_0775_, _0774_, _1470_);
    or _2327_(_0090_, _0775_, _0766_);
    and _2328_(_0776_, _1471_, packet_out[55]);
    and _2329_(_0777_, _1473_, packet_buffer_3[55]);
    and _2330_(_0778_, _1476_, packet_buffer_2[55]);
    or _2331_(_0779_, _0778_, _0777_);
    and _2332_(_0780_, _1479_, packet_buffer_1[55]);
    and _2333_(_0781_, _1481_, packet_buffer_0[55]);
    or _2334_(_0782_, _0781_, _0780_);
    or _2335_(_0783_, _0782_, _0779_);
    and _2336_(_0784_, _0783_, _1487_);
    and _2337_(_0785_, _0784_, _1470_);
    or _2338_(_0091_, _0785_, _0776_);
    and _2339_(_0786_, _1471_, packet_out[56]);
    and _2340_(_0787_, _1473_, packet_buffer_3[56]);
    and _2341_(_0788_, _1476_, packet_buffer_2[56]);
    or _2342_(_0789_, _0788_, _0787_);
    and _2343_(_0790_, _1479_, packet_buffer_1[56]);
    and _2344_(_0791_, _1481_, packet_buffer_0[56]);
    or _2345_(_0792_, _0791_, _0790_);
    or _2346_(_0793_, _0792_, _0789_);
    and _2347_(_0794_, _0793_, _1487_);
    and _2348_(_0795_, _0794_, _1470_);
    or _2349_(_0092_, _0795_, _0786_);
    and _2350_(_0796_, _1471_, packet_out[57]);
    and _2351_(_0797_, _1473_, packet_buffer_3[57]);
    and _2352_(_0798_, _1476_, packet_buffer_2[57]);
    or _2353_(_0799_, _0798_, _0797_);
    and _2354_(_0800_, _1479_, packet_buffer_1[57]);
    and _2355_(_0801_, _1481_, packet_buffer_0[57]);
    or _2356_(_0802_, _0801_, _0800_);
    or _2357_(_0803_, _0802_, _0799_);
    and _2358_(_0804_, _0803_, _1487_);
    and _2359_(_0805_, _0804_, _1470_);
    or _2360_(_0093_, _0805_, _0796_);
    and _2361_(_0806_, _1471_, packet_out[58]);
    and _2362_(_0807_, _1473_, packet_buffer_3[58]);
    and _2363_(_0808_, _1476_, packet_buffer_2[58]);
    or _2364_(_0809_, _0808_, _0807_);
    and _2365_(_0810_, _1479_, packet_buffer_1[58]);
    and _2366_(_0811_, _1481_, packet_buffer_0[58]);
    or _2367_(_0812_, _0811_, _0810_);
    or _2368_(_0813_, _0812_, _0809_);
    and _2369_(_0814_, _0813_, _1487_);
    and _2370_(_0815_, _0814_, _1470_);
    or _2371_(_0094_, _0815_, _0806_);
    and _2372_(_0816_, _1471_, packet_out[59]);
    and _2373_(_0817_, _1473_, packet_buffer_3[59]);
    and _2374_(_0818_, _1476_, packet_buffer_2[59]);
    or _2375_(_0819_, _0818_, _0817_);
    and _2376_(_0820_, _1479_, packet_buffer_1[59]);
    and _2377_(_0821_, _1481_, packet_buffer_0[59]);
    or _2378_(_0822_, _0821_, _0820_);
    or _2379_(_0823_, _0822_, _0819_);
    and _2380_(_0824_, _0823_, _1487_);
    and _2381_(_0825_, _0824_, _1470_);
    or _2382_(_0095_, _0825_, _0816_);
    and _2383_(_0826_, _1471_, packet_out[60]);
    and _2384_(_0827_, _1473_, packet_buffer_3[60]);
    and _2385_(_0828_, _1476_, packet_buffer_2[60]);
    or _2386_(_0829_, _0828_, _0827_);
    and _2387_(_0830_, _1479_, packet_buffer_1[60]);
    and _2388_(_0831_, _1481_, packet_buffer_0[60]);
    or _2389_(_0832_, _0831_, _0830_);
    or _2390_(_0833_, _0832_, _0829_);
    and _2391_(_0834_, _0833_, _1487_);
    and _2392_(_0835_, _0834_, _1470_);
    or _2393_(_0096_, _0835_, _0826_);
    and _2394_(_0836_, _1471_, packet_out[61]);
    and _2395_(_0837_, _1473_, packet_buffer_3[61]);
    and _2396_(_0838_, _1476_, packet_buffer_2[61]);
    or _2397_(_0839_, _0838_, _0837_);
    and _2398_(_0840_, _1479_, packet_buffer_1[61]);
    and _2399_(_0841_, _1481_, packet_buffer_0[61]);
    or _2400_(_0842_, _0841_, _0840_);
    or _2401_(_0843_, _0842_, _0839_);
    and _2402_(_0844_, _0843_, _1487_);
    and _2403_(_0845_, _0844_, _1470_);
    or _2404_(_0097_, _0845_, _0836_);
    and _2405_(_0846_, _1471_, packet_out[62]);
    and _2406_(_0847_, _1473_, packet_buffer_3[62]);
    and _2407_(_0848_, _1476_, packet_buffer_2[62]);
    or _2408_(_0849_, _0848_, _0847_);
    and _2409_(_0850_, _1479_, packet_buffer_1[62]);
    and _2410_(_0851_, _1481_, packet_buffer_0[62]);
    or _2411_(_0852_, _0851_, _0850_);
    or _2412_(_0853_, _0852_, _0849_);
    and _2413_(_0854_, _0853_, _1487_);
    and _2414_(_0855_, _0854_, _1470_);
    or _2415_(_0098_, _0855_, _0846_);
    and _2416_(_0856_, _1471_, packet_out[63]);
    and _2417_(_0857_, _1473_, packet_buffer_3[63]);
    and _2418_(_0858_, _1476_, packet_buffer_2[63]);
    or _2419_(_0859_, _0858_, _0857_);
    and _2420_(_0860_, _1479_, packet_buffer_1[63]);
    and _2421_(_0861_, _1481_, packet_buffer_0[63]);
    or _2422_(_0862_, _0861_, _0860_);
    or _2423_(_0863_, _0862_, _0859_);
    and _2424_(_0864_, _0863_, _1487_);
    and _2425_(_0865_, _0864_, _1470_);
    or _2426_(_0099_, _0865_, _0856_);
    not _2427_(_0866_, buffer_tail[1]);
    and _2428_(_0867_, _0866_, buffer_tail[0]);
    and _2429_(_0868_, _0867_, _1381_);
    not _2430_(_0869_, _0868_);
    and _2431_(_0870_, _0869_, packet_buffer_1[0]);
    and _2432_(_0871_, _0868_, packet_in[0]);
    or _2433_(_0100_, _0871_, _0870_);
    and _2434_(_0872_, _0869_, packet_buffer_1[1]);
    and _2435_(_0873_, _0868_, packet_in[1]);
    or _2436_(_0101_, _0873_, _0872_);
    and _2437_(_0874_, _0869_, packet_buffer_1[2]);
    and _2438_(_0875_, _0868_, packet_in[2]);
    or _2439_(_0102_, _0875_, _0874_);
    and _2440_(_0876_, _0869_, packet_buffer_1[3]);
    and _2441_(_0877_, _0868_, packet_in[3]);
    or _2442_(_0103_, _0877_, _0876_);
    and _2443_(_0878_, _0869_, packet_buffer_1[4]);
    and _2444_(_0879_, _0868_, packet_in[4]);
    or _2445_(_0104_, _0879_, _0878_);
    and _2446_(_0880_, _0869_, packet_buffer_1[5]);
    and _2447_(_0881_, _0868_, packet_in[5]);
    or _2448_(_0105_, _0881_, _0880_);
    and _2449_(_0882_, _0869_, packet_buffer_1[6]);
    and _2450_(_0883_, _0868_, packet_in[6]);
    or _2451_(_0106_, _0883_, _0882_);
    and _2452_(_0884_, _0869_, packet_buffer_1[7]);
    and _2453_(_0885_, _0868_, packet_in[7]);
    or _2454_(_0107_, _0885_, _0884_);
    and _2455_(_0886_, _0869_, packet_buffer_1[8]);
    and _2456_(_0887_, _0868_, packet_in[8]);
    or _2457_(_0108_, _0887_, _0886_);
    and _2458_(_0888_, _0869_, packet_buffer_1[9]);
    and _2459_(_0889_, _0868_, packet_in[9]);
    or _2460_(_0109_, _0889_, _0888_);
    and _2461_(_0890_, _0869_, packet_buffer_1[10]);
    and _2462_(_0891_, _0868_, packet_in[10]);
    or _2463_(_0110_, _0891_, _0890_);
    and _2464_(_0892_, _0869_, packet_buffer_1[11]);
    and _2465_(_0893_, _0868_, packet_in[11]);
    or _2466_(_0111_, _0893_, _0892_);
    and _2467_(_0894_, _0869_, packet_buffer_1[12]);
    and _2468_(_0895_, _0868_, packet_in[12]);
    or _2469_(_0112_, _0895_, _0894_);
    and _2470_(_0896_, _0869_, packet_buffer_1[13]);
    and _2471_(_0897_, _0868_, packet_in[13]);
    or _2472_(_0113_, _0897_, _0896_);
    and _2473_(_0898_, _0869_, packet_buffer_1[14]);
    and _2474_(_0899_, _0868_, packet_in[14]);
    or _2475_(_0114_, _0899_, _0898_);
    and _2476_(_0900_, _0869_, packet_buffer_1[15]);
    and _2477_(_0901_, _0868_, packet_in[15]);
    or _2478_(_0115_, _0901_, _0900_);
    and _2479_(_0902_, _0869_, packet_buffer_1[16]);
    and _2480_(_0903_, _0868_, packet_in[16]);
    or _2481_(_0116_, _0903_, _0902_);
    and _2482_(_0904_, _0869_, packet_buffer_1[17]);
    and _2483_(_0905_, _0868_, packet_in[17]);
    or _2484_(_0117_, _0905_, _0904_);
    and _2485_(_0906_, _0869_, packet_buffer_1[18]);
    and _2486_(_0907_, _0868_, packet_in[18]);
    or _2487_(_0118_, _0907_, _0906_);
    and _2488_(_0908_, _0869_, packet_buffer_1[19]);
    and _2489_(_0909_, _0868_, packet_in[19]);
    or _2490_(_0119_, _0909_, _0908_);
    and _2491_(_0910_, _0869_, packet_buffer_1[20]);
    and _2492_(_0911_, _0868_, packet_in[20]);
    or _2493_(_0120_, _0911_, _0910_);
    and _2494_(_0912_, _0869_, packet_buffer_1[21]);
    and _2495_(_0913_, _0868_, packet_in[21]);
    or _2496_(_0121_, _0913_, _0912_);
    and _2497_(_0914_, _0869_, packet_buffer_1[22]);
    and _2498_(_0915_, _0868_, packet_in[22]);
    or _2499_(_0122_, _0915_, _0914_);
    and _2500_(_0916_, _0869_, packet_buffer_1[23]);
    and _2501_(_0917_, _0868_, packet_in[23]);
    or _2502_(_0123_, _0917_, _0916_);
    and _2503_(_0918_, _0869_, packet_buffer_1[24]);
    and _2504_(_0919_, _0868_, packet_in[24]);
    or _2505_(_0124_, _0919_, _0918_);
    and _2506_(_0920_, _0869_, packet_buffer_1[25]);
    and _2507_(_0921_, _0868_, packet_in[25]);
    or _2508_(_0125_, _0921_, _0920_);
    and _2509_(_0922_, _0869_, packet_buffer_1[26]);
    and _2510_(_0923_, _0868_, packet_in[26]);
    or _2511_(_0126_, _0923_, _0922_);
    and _2512_(_0924_, _0869_, packet_buffer_1[27]);
    and _2513_(_0925_, _0868_, packet_in[27]);
    or _2514_(_0127_, _0925_, _0924_);
    and _2515_(_0926_, _0869_, packet_buffer_1[28]);
    and _2516_(_0927_, _0868_, packet_in[28]);
    or _2517_(_0128_, _0927_, _0926_);
    and _2518_(_0928_, _0869_, packet_buffer_1[29]);
    and _2519_(_0929_, _0868_, packet_in[29]);
    or _2520_(_0129_, _0929_, _0928_);
    and _2521_(_0930_, _0869_, packet_buffer_1[30]);
    and _2522_(_0931_, _0868_, packet_in[30]);
    or _2523_(_0130_, _0931_, _0930_);
    and _2524_(_0932_, _0869_, packet_buffer_1[31]);
    and _2525_(_0933_, _0868_, packet_in[31]);
    or _2526_(_0131_, _0933_, _0932_);
    and _2527_(_0934_, _0869_, packet_buffer_1[32]);
    and _2528_(_0935_, _0868_, packet_in[32]);
    or _2529_(_0132_, _0935_, _0934_);
    and _2530_(_0936_, _0869_, packet_buffer_1[33]);
    and _2531_(_0937_, _0868_, packet_in[33]);
    or _2532_(_0133_, _0937_, _0936_);
    and _2533_(_0938_, _0869_, packet_buffer_1[34]);
    and _2534_(_0939_, _0868_, packet_in[34]);
    or _2535_(_0134_, _0939_, _0938_);
    and _2536_(_0940_, _0869_, packet_buffer_1[35]);
    and _2537_(_0941_, _0868_, packet_in[35]);
    or _2538_(_0135_, _0941_, _0940_);
    and _2539_(_0942_, _0869_, packet_buffer_1[36]);
    and _2540_(_0943_, _0868_, packet_in[36]);
    or _2541_(_0136_, _0943_, _0942_);
    and _2542_(_0944_, _0869_, packet_buffer_1[37]);
    and _2543_(_0945_, _0868_, packet_in[37]);
    or _2544_(_0137_, _0945_, _0944_);
    and _2545_(_0946_, _0869_, packet_buffer_1[38]);
    and _2546_(_0947_, _0868_, packet_in[38]);
    or _2547_(_0138_, _0947_, _0946_);
    and _2548_(_0948_, _0869_, packet_buffer_1[39]);
    and _2549_(_0949_, _0868_, packet_in[39]);
    or _2550_(_0139_, _0949_, _0948_);
    and _2551_(_0950_, _0869_, packet_buffer_1[40]);
    and _2552_(_0951_, _0868_, packet_in[40]);
    or _2553_(_0140_, _0951_, _0950_);
    and _2554_(_0952_, _0869_, packet_buffer_1[41]);
    and _2555_(_0953_, _0868_, packet_in[41]);
    or _2556_(_0141_, _0953_, _0952_);
    and _2557_(_0954_, _0869_, packet_buffer_1[42]);
    and _2558_(_0955_, _0868_, packet_in[42]);
    or _2559_(_0142_, _0955_, _0954_);
    and _2560_(_0956_, _0869_, packet_buffer_1[43]);
    and _2561_(_0957_, _0868_, packet_in[43]);
    or _2562_(_0143_, _0957_, _0956_);
    and _2563_(_0958_, _0869_, packet_buffer_1[44]);
    and _2564_(_0959_, _0868_, packet_in[44]);
    or _2565_(_0144_, _0959_, _0958_);
    and _2566_(_0960_, _0869_, packet_buffer_1[45]);
    and _2567_(_0961_, _0868_, packet_in[45]);
    or _2568_(_0145_, _0961_, _0960_);
    and _2569_(_0962_, _0869_, packet_buffer_1[46]);
    and _2570_(_0963_, _0868_, packet_in[46]);
    or _2571_(_0146_, _0963_, _0962_);
    and _2572_(_0964_, _0869_, packet_buffer_1[47]);
    and _2573_(_0965_, _0868_, packet_in[47]);
    or _2574_(_0147_, _0965_, _0964_);
    and _2575_(_0966_, _0869_, packet_buffer_1[48]);
    and _2576_(_0967_, _0868_, packet_in[48]);
    or _2577_(_0148_, _0967_, _0966_);
    and _2578_(_0968_, _0869_, packet_buffer_1[49]);
    and _2579_(_0969_, _0868_, packet_in[49]);
    or _2580_(_0149_, _0969_, _0968_);
    and _2581_(_0970_, _0869_, packet_buffer_1[50]);
    and _2582_(_0971_, _0868_, packet_in[50]);
    or _2583_(_0150_, _0971_, _0970_);
    and _2584_(_0972_, _0869_, packet_buffer_1[51]);
    and _2585_(_0973_, _0868_, packet_in[51]);
    or _2586_(_0151_, _0973_, _0972_);
    and _2587_(_0974_, _0869_, packet_buffer_1[52]);
    and _2588_(_0975_, _0868_, packet_in[52]);
    or _2589_(_0152_, _0975_, _0974_);
    and _2590_(_0976_, _0869_, packet_buffer_1[53]);
    and _2591_(_0977_, _0868_, packet_in[53]);
    or _2592_(_0153_, _0977_, _0976_);
    and _2593_(_0978_, _0869_, packet_buffer_1[54]);
    and _2594_(_0979_, _0868_, packet_in[54]);
    or _2595_(_0154_, _0979_, _0978_);
    and _2596_(_0980_, _0869_, packet_buffer_1[55]);
    and _2597_(_0981_, _0868_, packet_in[55]);
    or _2598_(_0155_, _0981_, _0980_);
    and _2599_(_0982_, _0869_, packet_buffer_1[56]);
    and _2600_(_0983_, _0868_, packet_in[56]);
    or _2601_(_0156_, _0983_, _0982_);
    and _2602_(_0984_, _0869_, packet_buffer_1[57]);
    and _2603_(_0985_, _0868_, packet_in[57]);
    or _2604_(_0157_, _0985_, _0984_);
    and _2605_(_0986_, _0869_, packet_buffer_1[58]);
    and _2606_(_0987_, _0868_, packet_in[58]);
    or _2607_(_0158_, _0987_, _0986_);
    and _2608_(_0988_, _0869_, packet_buffer_1[59]);
    and _2609_(_0989_, _0868_, packet_in[59]);
    or _2610_(_0159_, _0989_, _0988_);
    and _2611_(_0990_, _0869_, packet_buffer_1[60]);
    and _2612_(_0991_, _0868_, packet_in[60]);
    or _2613_(_0160_, _0991_, _0990_);
    and _2614_(_0992_, _0869_, packet_buffer_1[61]);
    and _2615_(_0993_, _0868_, packet_in[61]);
    or _2616_(_0161_, _0993_, _0992_);
    and _2617_(_0994_, _0869_, packet_buffer_1[62]);
    and _2618_(_0995_, _0868_, packet_in[62]);
    or _2619_(_0162_, _0995_, _0994_);
    and _2620_(_0996_, _0869_, packet_buffer_1[63]);
    and _2621_(_0997_, _0868_, packet_in[63]);
    or _2622_(_0163_, _0997_, _0996_);
    nor _2623_(_0998_, _1450_, _1410_);
    and _2624_(_0999_, _0998_, packet_ready);
    and _2625_(_1000_, _1409_, _1377_);
    or _2626_(_0164_, _1000_, _0999_);
    nor _2627_(_1001_, buffer_tail[1], buffer_tail[0]);
    and _2628_(_1002_, _1001_, _1381_);
    not _2629_(_1003_, _1002_);
    and _2630_(_1004_, _1003_, packet_buffer_0[0]);
    and _2631_(_1005_, _1002_, packet_in[0]);
    or _2632_(_0166_, _1005_, _1004_);
    and _2633_(_1006_, _1003_, packet_buffer_0[1]);
    and _2634_(_1007_, _1002_, packet_in[1]);
    or _2635_(_0167_, _1007_, _1006_);
    and _2636_(_1008_, _1003_, packet_buffer_0[2]);
    and _2637_(_1009_, _1002_, packet_in[2]);
    or _2638_(_0168_, _1009_, _1008_);
    and _2639_(_1010_, _1003_, packet_buffer_0[3]);
    and _2640_(_1011_, _1002_, packet_in[3]);
    or _2641_(_0169_, _1011_, _1010_);
    and _2642_(_1012_, _1003_, packet_buffer_0[4]);
    and _2643_(_1013_, _1002_, packet_in[4]);
    or _2644_(_0170_, _1013_, _1012_);
    and _2645_(_1014_, _1003_, packet_buffer_0[5]);
    and _2646_(_1015_, _1002_, packet_in[5]);
    or _2647_(_0171_, _1015_, _1014_);
    and _2648_(_1016_, _1003_, packet_buffer_0[6]);
    and _2649_(_1017_, _1002_, packet_in[6]);
    or _2650_(_0172_, _1017_, _1016_);
    and _2651_(_1018_, _1003_, packet_buffer_0[7]);
    and _2652_(_1019_, _1002_, packet_in[7]);
    or _2653_(_0173_, _1019_, _1018_);
    and _2654_(_1020_, _1003_, packet_buffer_0[8]);
    and _2655_(_1021_, _1002_, packet_in[8]);
    or _2656_(_0174_, _1021_, _1020_);
    and _2657_(_1022_, _1003_, packet_buffer_0[9]);
    and _2658_(_1023_, _1002_, packet_in[9]);
    or _2659_(_0175_, _1023_, _1022_);
    and _2660_(_1024_, _1003_, packet_buffer_0[10]);
    and _2661_(_1025_, _1002_, packet_in[10]);
    or _2662_(_0176_, _1025_, _1024_);
    and _2663_(_1026_, _1003_, packet_buffer_0[11]);
    and _2664_(_1027_, _1002_, packet_in[11]);
    or _2665_(_0177_, _1027_, _1026_);
    and _2666_(_1028_, _1003_, packet_buffer_0[12]);
    and _2667_(_1029_, _1002_, packet_in[12]);
    or _2668_(_0178_, _1029_, _1028_);
    and _2669_(_1030_, _1003_, packet_buffer_0[13]);
    and _2670_(_1031_, _1002_, packet_in[13]);
    or _2671_(_0179_, _1031_, _1030_);
    and _2672_(_1032_, _1003_, packet_buffer_0[14]);
    and _2673_(_1033_, _1002_, packet_in[14]);
    or _2674_(_0180_, _1033_, _1032_);
    and _2675_(_1034_, _1003_, packet_buffer_0[15]);
    and _2676_(_1035_, _1002_, packet_in[15]);
    or _2677_(_0181_, _1035_, _1034_);
    and _2678_(_1036_, _1003_, packet_buffer_0[16]);
    and _2679_(_1037_, _1002_, packet_in[16]);
    or _2680_(_0182_, _1037_, _1036_);
    and _2681_(_1038_, _1003_, packet_buffer_0[17]);
    and _2682_(_1039_, _1002_, packet_in[17]);
    or _2683_(_0183_, _1039_, _1038_);
    and _2684_(_1040_, _1003_, packet_buffer_0[18]);
    and _2685_(_1041_, _1002_, packet_in[18]);
    or _2686_(_0184_, _1041_, _1040_);
    and _2687_(_1042_, _1003_, packet_buffer_0[19]);
    and _2688_(_1043_, _1002_, packet_in[19]);
    or _2689_(_0185_, _1043_, _1042_);
    and _2690_(_1044_, _1003_, packet_buffer_0[20]);
    and _2691_(_1045_, _1002_, packet_in[20]);
    or _2692_(_0186_, _1045_, _1044_);
    and _2693_(_1046_, _1003_, packet_buffer_0[21]);
    and _2694_(_1047_, _1002_, packet_in[21]);
    or _2695_(_0187_, _1047_, _1046_);
    and _2696_(_1048_, _1003_, packet_buffer_0[22]);
    and _2697_(_1049_, _1002_, packet_in[22]);
    or _2698_(_0188_, _1049_, _1048_);
    and _2699_(_1050_, _1003_, packet_buffer_0[23]);
    and _2700_(_1051_, _1002_, packet_in[23]);
    or _2701_(_0189_, _1051_, _1050_);
    and _2702_(_1052_, _1003_, packet_buffer_0[24]);
    and _2703_(_1053_, _1002_, packet_in[24]);
    or _2704_(_0190_, _1053_, _1052_);
    and _2705_(_1054_, _1003_, packet_buffer_0[25]);
    and _2706_(_1055_, _1002_, packet_in[25]);
    or _2707_(_0191_, _1055_, _1054_);
    and _2708_(_1056_, _1003_, packet_buffer_0[26]);
    and _2709_(_1057_, _1002_, packet_in[26]);
    or _2710_(_0192_, _1057_, _1056_);
    and _2711_(_1058_, _1003_, packet_buffer_0[27]);
    and _2712_(_1059_, _1002_, packet_in[27]);
    or _2713_(_0193_, _1059_, _1058_);
    and _2714_(_1060_, _1003_, packet_buffer_0[28]);
    and _2715_(_1061_, _1002_, packet_in[28]);
    or _2716_(_0194_, _1061_, _1060_);
    and _2717_(_1062_, _1003_, packet_buffer_0[29]);
    and _2718_(_1063_, _1002_, packet_in[29]);
    or _2719_(_0195_, _1063_, _1062_);
    and _2720_(_1064_, _1003_, packet_buffer_0[30]);
    and _2721_(_1065_, _1002_, packet_in[30]);
    or _2722_(_0196_, _1065_, _1064_);
    and _2723_(_1066_, _1003_, packet_buffer_0[31]);
    and _2724_(_1067_, _1002_, packet_in[31]);
    or _2725_(_0197_, _1067_, _1066_);
    and _2726_(_1068_, _1003_, packet_buffer_0[32]);
    and _2727_(_1069_, _1002_, packet_in[32]);
    or _2728_(_0198_, _1069_, _1068_);
    and _2729_(_1070_, _1003_, packet_buffer_0[33]);
    and _2730_(_1071_, _1002_, packet_in[33]);
    or _2731_(_0199_, _1071_, _1070_);
    and _2732_(_1072_, _1003_, packet_buffer_0[34]);
    and _2733_(_1073_, _1002_, packet_in[34]);
    or _2734_(_0200_, _1073_, _1072_);
    and _2735_(_1074_, _1003_, packet_buffer_0[35]);
    and _2736_(_1075_, _1002_, packet_in[35]);
    or _2737_(_0201_, _1075_, _1074_);
    and _2738_(_1076_, _1003_, packet_buffer_0[36]);
    and _2739_(_1077_, _1002_, packet_in[36]);
    or _2740_(_0202_, _1077_, _1076_);
    and _2741_(_1078_, _1003_, packet_buffer_0[37]);
    and _2742_(_1079_, _1002_, packet_in[37]);
    or _2743_(_0203_, _1079_, _1078_);
    and _2744_(_1080_, _1003_, packet_buffer_0[38]);
    and _2745_(_1081_, _1002_, packet_in[38]);
    or _2746_(_0204_, _1081_, _1080_);
    and _2747_(_1082_, _1003_, packet_buffer_0[39]);
    and _2748_(_1083_, _1002_, packet_in[39]);
    or _2749_(_0205_, _1083_, _1082_);
    and _2750_(_1084_, _1003_, packet_buffer_0[40]);
    and _2751_(_1085_, _1002_, packet_in[40]);
    or _2752_(_0206_, _1085_, _1084_);
    and _2753_(_1086_, _1003_, packet_buffer_0[41]);
    and _2754_(_1087_, _1002_, packet_in[41]);
    or _2755_(_0207_, _1087_, _1086_);
    and _2756_(_1088_, _1003_, packet_buffer_0[42]);
    and _2757_(_1089_, _1002_, packet_in[42]);
    or _2758_(_0208_, _1089_, _1088_);
    and _2759_(_1090_, _1003_, packet_buffer_0[43]);
    and _2760_(_1091_, _1002_, packet_in[43]);
    or _2761_(_0209_, _1091_, _1090_);
    and _2762_(_1092_, _1003_, packet_buffer_0[44]);
    and _2763_(_1093_, _1002_, packet_in[44]);
    or _2764_(_0210_, _1093_, _1092_);
    and _2765_(_1094_, _1003_, packet_buffer_0[45]);
    and _2766_(_1095_, _1002_, packet_in[45]);
    or _2767_(_0211_, _1095_, _1094_);
    and _2768_(_1096_, _1003_, packet_buffer_0[46]);
    and _2769_(_1097_, _1002_, packet_in[46]);
    or _2770_(_0212_, _1097_, _1096_);
    and _2771_(_1098_, _1003_, packet_buffer_0[47]);
    and _2772_(_1099_, _1002_, packet_in[47]);
    or _2773_(_0213_, _1099_, _1098_);
    and _2774_(_1100_, _1003_, packet_buffer_0[48]);
    and _2775_(_1101_, _1002_, packet_in[48]);
    or _2776_(_0214_, _1101_, _1100_);
    and _2777_(_1102_, _1003_, packet_buffer_0[49]);
    and _2778_(_1103_, _1002_, packet_in[49]);
    or _2779_(_0215_, _1103_, _1102_);
    and _2780_(_1104_, _1003_, packet_buffer_0[50]);
    and _2781_(_1105_, _1002_, packet_in[50]);
    or _2782_(_0216_, _1105_, _1104_);
    and _2783_(_1106_, _1003_, packet_buffer_0[51]);
    and _2784_(_1107_, _1002_, packet_in[51]);
    or _2785_(_0217_, _1107_, _1106_);
    and _2786_(_1108_, _1003_, packet_buffer_0[52]);
    and _2787_(_1109_, _1002_, packet_in[52]);
    or _2788_(_0218_, _1109_, _1108_);
    and _2789_(_1110_, _1003_, packet_buffer_0[53]);
    and _2790_(_1111_, _1002_, packet_in[53]);
    or _2791_(_0219_, _1111_, _1110_);
    and _2792_(_1112_, _1003_, packet_buffer_0[54]);
    and _2793_(_1113_, _1002_, packet_in[54]);
    or _2794_(_0220_, _1113_, _1112_);
    and _2795_(_1114_, _1003_, packet_buffer_0[55]);
    and _2796_(_1115_, _1002_, packet_in[55]);
    or _2797_(_0221_, _1115_, _1114_);
    and _2798_(_1116_, _1003_, packet_buffer_0[56]);
    and _2799_(_1117_, _1002_, packet_in[56]);
    or _2800_(_0222_, _1117_, _1116_);
    and _2801_(_1118_, _1003_, packet_buffer_0[57]);
    and _2802_(_1119_, _1002_, packet_in[57]);
    or _2803_(_0223_, _1119_, _1118_);
    and _2804_(_1120_, _1003_, packet_buffer_0[58]);
    and _2805_(_1121_, _1002_, packet_in[58]);
    or _2806_(_0224_, _1121_, _1120_);
    and _2807_(_1122_, _1003_, packet_buffer_0[59]);
    and _2808_(_1123_, _1002_, packet_in[59]);
    or _2809_(_0225_, _1123_, _1122_);
    and _2810_(_1124_, _1003_, packet_buffer_0[60]);
    and _2811_(_1125_, _1002_, packet_in[60]);
    or _2812_(_0226_, _1125_, _1124_);
    and _2813_(_1126_, _1003_, packet_buffer_0[61]);
    and _2814_(_1127_, _1002_, packet_in[61]);
    or _2815_(_0227_, _1127_, _1126_);
    and _2816_(_1128_, _1003_, packet_buffer_0[62]);
    and _2817_(_1129_, _1002_, packet_in[62]);
    or _2818_(_0228_, _1129_, _1128_);
    and _2819_(_1130_, _1003_, packet_buffer_0[63]);
    and _2820_(_1131_, _1002_, packet_in[63]);
    or _2821_(_0229_, _1131_, _1130_);
    nor _2822_(_1132_, _0866_, buffer_tail[0]);
    and _2823_(_1133_, _1132_, _1381_);
    not _2824_(_1134_, _1133_);
    and _2825_(_1135_, _1134_, packet_buffer_2[0]);
    and _2826_(_1136_, _1133_, packet_in[0]);
    or _2827_(_0230_, _1136_, _1135_);
    and _2828_(_1137_, _1134_, packet_buffer_2[1]);
    and _2829_(_1138_, _1133_, packet_in[1]);
    or _2830_(_0231_, _1138_, _1137_);
    and _2831_(_1139_, _1134_, packet_buffer_2[2]);
    and _2832_(_1140_, _1133_, packet_in[2]);
    or _2833_(_0232_, _1140_, _1139_);
    and _2834_(_1141_, _1134_, packet_buffer_2[3]);
    and _2835_(_1142_, _1133_, packet_in[3]);
    or _2836_(_0233_, _1142_, _1141_);
    and _2837_(_1143_, _1134_, packet_buffer_2[4]);
    and _2838_(_1144_, _1133_, packet_in[4]);
    or _2839_(_0234_, _1144_, _1143_);
    and _2840_(_1145_, _1134_, packet_buffer_2[5]);
    and _2841_(_1146_, _1133_, packet_in[5]);
    or _2842_(_0235_, _1146_, _1145_);
    and _2843_(_1147_, _1134_, packet_buffer_2[6]);
    and _2844_(_1148_, _1133_, packet_in[6]);
    or _2845_(_0236_, _1148_, _1147_);
    and _2846_(_1149_, _1134_, packet_buffer_2[7]);
    and _2847_(_1150_, _1133_, packet_in[7]);
    or _2848_(_0237_, _1150_, _1149_);
    and _2849_(_1151_, _1134_, packet_buffer_2[8]);
    and _2850_(_1152_, _1133_, packet_in[8]);
    or _2851_(_0238_, _1152_, _1151_);
    and _2852_(_1153_, _1134_, packet_buffer_2[9]);
    and _2853_(_1154_, _1133_, packet_in[9]);
    or _2854_(_0239_, _1154_, _1153_);
    and _2855_(_1155_, _1134_, packet_buffer_2[10]);
    and _2856_(_1156_, _1133_, packet_in[10]);
    or _2857_(_0240_, _1156_, _1155_);
    and _2858_(_1157_, _1134_, packet_buffer_2[11]);
    and _2859_(_1158_, _1133_, packet_in[11]);
    or _2860_(_0241_, _1158_, _1157_);
    and _2861_(_1159_, _1134_, packet_buffer_2[12]);
    and _2862_(_1160_, _1133_, packet_in[12]);
    or _2863_(_0242_, _1160_, _1159_);
    and _2864_(_1161_, _1134_, packet_buffer_2[13]);
    and _2865_(_1162_, _1133_, packet_in[13]);
    or _2866_(_0243_, _1162_, _1161_);
    and _2867_(_1163_, _1134_, packet_buffer_2[14]);
    and _2868_(_1164_, _1133_, packet_in[14]);
    or _2869_(_0244_, _1164_, _1163_);
    and _2870_(_1165_, _1134_, packet_buffer_2[15]);
    and _2871_(_1166_, _1133_, packet_in[15]);
    or _2872_(_0245_, _1166_, _1165_);
    and _2873_(_1167_, _1134_, packet_buffer_2[16]);
    and _2874_(_1168_, _1133_, packet_in[16]);
    or _2875_(_0246_, _1168_, _1167_);
    and _2876_(_1169_, _1134_, packet_buffer_2[17]);
    and _2877_(_1170_, _1133_, packet_in[17]);
    or _2878_(_0247_, _1170_, _1169_);
    and _2879_(_1171_, _1134_, packet_buffer_2[18]);
    and _2880_(_1172_, _1133_, packet_in[18]);
    or _2881_(_0248_, _1172_, _1171_);
    and _2882_(_1173_, _1134_, packet_buffer_2[19]);
    and _2883_(_1174_, _1133_, packet_in[19]);
    or _2884_(_0249_, _1174_, _1173_);
    and _2885_(_1175_, _1134_, packet_buffer_2[20]);
    and _2886_(_1176_, _1133_, packet_in[20]);
    or _2887_(_0250_, _1176_, _1175_);
    and _2888_(_1177_, _1134_, packet_buffer_2[21]);
    and _2889_(_1178_, _1133_, packet_in[21]);
    or _2890_(_0251_, _1178_, _1177_);
    and _2891_(_1179_, _1134_, packet_buffer_2[22]);
    and _2892_(_1180_, _1133_, packet_in[22]);
    or _2893_(_0252_, _1180_, _1179_);
    and _2894_(_1181_, _1134_, packet_buffer_2[23]);
    and _2895_(_1182_, _1133_, packet_in[23]);
    or _2896_(_0253_, _1182_, _1181_);
    and _2897_(_1183_, _1134_, packet_buffer_2[24]);
    and _2898_(_1184_, _1133_, packet_in[24]);
    or _2899_(_0254_, _1184_, _1183_);
    and _2900_(_1185_, _1134_, packet_buffer_2[25]);
    and _2901_(_1186_, _1133_, packet_in[25]);
    or _2902_(_0255_, _1186_, _1185_);
    and _2903_(_1187_, _1134_, packet_buffer_2[26]);
    and _2904_(_1188_, _1133_, packet_in[26]);
    or _2905_(_0256_, _1188_, _1187_);
    and _2906_(_1189_, _1134_, packet_buffer_2[27]);
    and _2907_(_1190_, _1133_, packet_in[27]);
    or _2908_(_0257_, _1190_, _1189_);
    and _2909_(_1191_, _1134_, packet_buffer_2[28]);
    and _2910_(_1192_, _1133_, packet_in[28]);
    or _2911_(_0258_, _1192_, _1191_);
    and _2912_(_1193_, _1134_, packet_buffer_2[29]);
    and _2913_(_1194_, _1133_, packet_in[29]);
    or _2914_(_0259_, _1194_, _1193_);
    and _2915_(_1195_, _1134_, packet_buffer_2[30]);
    and _2916_(_1196_, _1133_, packet_in[30]);
    or _2917_(_0260_, _1196_, _1195_);
    and _2918_(_1197_, _1134_, packet_buffer_2[31]);
    and _2919_(_1198_, _1133_, packet_in[31]);
    or _2920_(_0261_, _1198_, _1197_);
    and _2921_(_1199_, _1134_, packet_buffer_2[32]);
    and _2922_(_1200_, _1133_, packet_in[32]);
    or _2923_(_0262_, _1200_, _1199_);
    and _2924_(_1201_, _1134_, packet_buffer_2[33]);
    and _2925_(_1202_, _1133_, packet_in[33]);
    or _2926_(_0263_, _1202_, _1201_);
    and _2927_(_1203_, _1134_, packet_buffer_2[34]);
    and _2928_(_1204_, _1133_, packet_in[34]);
    or _2929_(_0264_, _1204_, _1203_);
    and _2930_(_1205_, _1134_, packet_buffer_2[35]);
    and _2931_(_1206_, _1133_, packet_in[35]);
    or _2932_(_0265_, _1206_, _1205_);
    and _2933_(_1207_, _1134_, packet_buffer_2[36]);
    and _2934_(_1208_, _1133_, packet_in[36]);
    or _2935_(_0266_, _1208_, _1207_);
    and _2936_(_1209_, _1134_, packet_buffer_2[37]);
    and _2937_(_1210_, _1133_, packet_in[37]);
    or _2938_(_0267_, _1210_, _1209_);
    and _2939_(_1211_, _1134_, packet_buffer_2[38]);
    and _2940_(_1212_, _1133_, packet_in[38]);
    or _2941_(_0268_, _1212_, _1211_);
    and _2942_(_1213_, _1134_, packet_buffer_2[39]);
    and _2943_(_1214_, _1133_, packet_in[39]);
    or _2944_(_0269_, _1214_, _1213_);
    and _2945_(_1215_, _1134_, packet_buffer_2[40]);
    and _2946_(_1216_, _1133_, packet_in[40]);
    or _2947_(_0270_, _1216_, _1215_);
    and _2948_(_1217_, _1134_, packet_buffer_2[41]);
    and _2949_(_1218_, _1133_, packet_in[41]);
    or _2950_(_0271_, _1218_, _1217_);
    and _2951_(_1219_, _1134_, packet_buffer_2[42]);
    and _2952_(_1220_, _1133_, packet_in[42]);
    or _2953_(_0272_, _1220_, _1219_);
    and _2954_(_1221_, _1134_, packet_buffer_2[43]);
    and _2955_(_1222_, _1133_, packet_in[43]);
    or _2956_(_0273_, _1222_, _1221_);
    and _2957_(_1223_, _1134_, packet_buffer_2[44]);
    and _2958_(_1224_, _1133_, packet_in[44]);
    or _2959_(_0274_, _1224_, _1223_);
    and _2960_(_1225_, _1134_, packet_buffer_2[45]);
    and _2961_(_1226_, _1133_, packet_in[45]);
    or _2962_(_0275_, _1226_, _1225_);
    and _2963_(_1227_, _1134_, packet_buffer_2[46]);
    and _2964_(_1228_, _1133_, packet_in[46]);
    or _2965_(_0276_, _1228_, _1227_);
    and _2966_(_1229_, _1134_, packet_buffer_2[47]);
    and _2967_(_1230_, _1133_, packet_in[47]);
    or _2968_(_0277_, _1230_, _1229_);
    and _2969_(_1231_, _1134_, packet_buffer_2[48]);
    and _2970_(_1232_, _1133_, packet_in[48]);
    or _2971_(_0278_, _1232_, _1231_);
    and _2972_(_1233_, _1134_, packet_buffer_2[49]);
    and _2973_(_1234_, _1133_, packet_in[49]);
    or _2974_(_0279_, _1234_, _1233_);
    and _2975_(_1235_, _1134_, packet_buffer_2[50]);
    and _2976_(_1236_, _1133_, packet_in[50]);
    or _2977_(_0280_, _1236_, _1235_);
    and _2978_(_1237_, _1134_, packet_buffer_2[51]);
    and _2979_(_1238_, _1133_, packet_in[51]);
    or _2980_(_0281_, _1238_, _1237_);
    and _2981_(_1239_, _1134_, packet_buffer_2[52]);
    and _2982_(_1240_, _1133_, packet_in[52]);
    or _2983_(_0282_, _1240_, _1239_);
    and _2984_(_1241_, _1134_, packet_buffer_2[53]);
    and _2985_(_1242_, _1133_, packet_in[53]);
    or _2986_(_0283_, _1242_, _1241_);
    and _2987_(_1243_, _1134_, packet_buffer_2[54]);
    and _2988_(_1244_, _1133_, packet_in[54]);
    or _2989_(_0284_, _1244_, _1243_);
    and _2990_(_1245_, _1134_, packet_buffer_2[55]);
    and _2991_(_1246_, _1133_, packet_in[55]);
    or _2992_(_0285_, _1246_, _1245_);
    and _2993_(_1247_, _1134_, packet_buffer_2[56]);
    and _2994_(_1248_, _1133_, packet_in[56]);
    or _2995_(_0286_, _1248_, _1247_);
    and _2996_(_1249_, _1134_, packet_buffer_2[57]);
    and _2997_(_1250_, _1133_, packet_in[57]);
    or _2998_(_0287_, _1250_, _1249_);
    and _2999_(_1251_, _1134_, packet_buffer_2[58]);
    and _3000_(_1252_, _1133_, packet_in[58]);
    or _3001_(_0288_, _1252_, _1251_);
    and _3002_(_1253_, _1134_, packet_buffer_2[59]);
    and _3003_(_1254_, _1133_, packet_in[59]);
    or _3004_(_0289_, _1254_, _1253_);
    and _3005_(_1255_, _1134_, packet_buffer_2[60]);
    and _3006_(_1256_, _1133_, packet_in[60]);
    or _3007_(_0290_, _1256_, _1255_);
    and _3008_(_1257_, _1134_, packet_buffer_2[61]);
    and _3009_(_1258_, _1133_, packet_in[61]);
    or _3010_(_0291_, _1258_, _1257_);
    and _3011_(_1259_, _1134_, packet_buffer_2[62]);
    and _3012_(_1260_, _1133_, packet_in[62]);
    or _3013_(_0292_, _1260_, _1259_);
    and _3014_(_1261_, _1134_, packet_buffer_2[63]);
    and _3015_(_1262_, _1133_, packet_in[63]);
    or _3016_(_0293_, _1262_, _1261_);
    and _3017_(_1263_, _1384_, packet_buffer_3[0]);
    and _3018_(_1264_, _1383_, packet_in[0]);
    or _3019_(_0294_, _1264_, _1263_);
    and _3020_(_1265_, _1384_, packet_buffer_3[1]);
    and _3021_(_1266_, _1383_, packet_in[1]);
    or _3022_(_0295_, _1266_, _1265_);
    and _3023_(_1267_, _1384_, packet_buffer_3[2]);
    and _3024_(_1268_, _1383_, packet_in[2]);
    or _3025_(_0296_, _1268_, _1267_);
    and _3026_(_1269_, _1384_, packet_buffer_3[3]);
    and _3027_(_1270_, _1383_, packet_in[3]);
    or _3028_(_0297_, _1270_, _1269_);
    and _3029_(_1271_, _1384_, packet_buffer_3[4]);
    and _3030_(_1272_, _1383_, packet_in[4]);
    or _3031_(_0298_, _1272_, _1271_);
    and _3032_(_1273_, _1384_, packet_buffer_3[5]);
    and _3033_(_1274_, _1383_, packet_in[5]);
    or _3034_(_0299_, _1274_, _1273_);
    and _3035_(_1275_, _1384_, packet_buffer_3[6]);
    and _3036_(_1276_, _1383_, packet_in[6]);
    or _3037_(_0300_, _1276_, _1275_);
    and _3038_(_1277_, _1384_, packet_buffer_3[7]);
    and _3039_(_1278_, _1383_, packet_in[7]);
    or _3040_(_0301_, _1278_, _1277_);
    and _3041_(_1279_, _1384_, packet_buffer_3[8]);
    and _3042_(_1280_, _1383_, packet_in[8]);
    or _3043_(_0302_, _1280_, _1279_);
    and _3044_(_1281_, _1384_, packet_buffer_3[9]);
    and _3045_(_1282_, _1383_, packet_in[9]);
    or _3046_(_0303_, _1282_, _1281_);
    and _3047_(_1283_, _1384_, packet_buffer_3[10]);
    and _3048_(_1284_, _1383_, packet_in[10]);
    or _3049_(_0304_, _1284_, _1283_);
    and _3050_(_1285_, _1384_, packet_buffer_3[11]);
    and _3051_(_1286_, _1383_, packet_in[11]);
    or _3052_(_0305_, _1286_, _1285_);
    and _3053_(_1287_, _1384_, packet_buffer_3[12]);
    and _3054_(_1288_, _1383_, packet_in[12]);
    or _3055_(_0306_, _1288_, _1287_);
    and _3056_(_1289_, _1384_, packet_buffer_3[13]);
    and _3057_(_1290_, _1383_, packet_in[13]);
    or _3058_(_0307_, _1290_, _1289_);
    and _3059_(_1291_, _1384_, packet_buffer_3[14]);
    and _3060_(_1292_, _1383_, packet_in[14]);
    or _3061_(_0308_, _1292_, _1291_);
    and _3062_(_1293_, _1384_, packet_buffer_3[15]);
    and _3063_(_1294_, _1383_, packet_in[15]);
    or _3064_(_0309_, _1294_, _1293_);
    and _3065_(_1295_, _1384_, packet_buffer_3[16]);
    and _3066_(_1296_, _1383_, packet_in[16]);
    or _3067_(_0310_, _1296_, _1295_);
    and _3068_(_1297_, _1384_, packet_buffer_3[17]);
    and _3069_(_1298_, _1383_, packet_in[17]);
    or _3070_(_0311_, _1298_, _1297_);
    and _3071_(_1299_, _1384_, packet_buffer_3[18]);
    and _3072_(_1300_, _1383_, packet_in[18]);
    or _3073_(_0312_, _1300_, _1299_);
    and _3074_(_1301_, _1384_, packet_buffer_3[19]);
    and _3075_(_1302_, _1383_, packet_in[19]);
    or _3076_(_0313_, _1302_, _1301_);
    and _3077_(_1303_, _1384_, packet_buffer_3[20]);
    and _3078_(_1304_, _1383_, packet_in[20]);
    or _3079_(_0314_, _1304_, _1303_);
    and _3080_(_1305_, _1384_, packet_buffer_3[21]);
    and _3081_(_1306_, _1383_, packet_in[21]);
    or _3082_(_0315_, _1306_, _1305_);
    and _3083_(_1307_, _1384_, packet_buffer_3[22]);
    and _3084_(_1308_, _1383_, packet_in[22]);
    or _3085_(_0316_, _1308_, _1307_);
    and _3086_(_1309_, _1384_, packet_buffer_3[23]);
    and _3087_(_1310_, _1383_, packet_in[23]);
    or _3088_(_0317_, _1310_, _1309_);
    and _3089_(_1311_, _1384_, packet_buffer_3[24]);
    and _3090_(_1312_, _1383_, packet_in[24]);
    or _3091_(_0318_, _1312_, _1311_);
    and _3092_(_1313_, _1384_, packet_buffer_3[25]);
    and _3093_(_1314_, _1383_, packet_in[25]);
    or _3094_(_0319_, _1314_, _1313_);
    and _3095_(_1315_, _1384_, packet_buffer_3[26]);
    and _3096_(_1316_, _1383_, packet_in[26]);
    or _3097_(_0320_, _1316_, _1315_);
    and _3098_(_1317_, _1384_, packet_buffer_3[27]);
    and _3099_(_1318_, _1383_, packet_in[27]);
    or _3100_(_0321_, _1318_, _1317_);
    and _3101_(_1319_, _1384_, packet_buffer_3[28]);
    and _3102_(_1320_, _1383_, packet_in[28]);
    or _3103_(_0322_, _1320_, _1319_);
    and _3104_(_1321_, _1384_, packet_buffer_3[29]);
    and _3105_(_1322_, _1383_, packet_in[29]);
    or _3106_(_0323_, _1322_, _1321_);
    and _3107_(_1323_, _1384_, packet_buffer_3[30]);
    and _3108_(_1324_, _1383_, packet_in[30]);
    or _3109_(_0324_, _1324_, _1323_);
    and _3110_(_1325_, _1384_, packet_buffer_3[31]);
    and _3111_(_1326_, _1383_, packet_in[31]);
    or _3112_(_0325_, _1326_, _1325_);
    and _3113_(_1327_, _1384_, packet_buffer_3[32]);
    and _3114_(_1328_, _1383_, packet_in[32]);
    or _3115_(_0326_, _1328_, _1327_);
    and _3116_(_1329_, _1384_, packet_buffer_3[33]);
    and _3117_(_1330_, _1383_, packet_in[33]);
    or _3118_(_0327_, _1330_, _1329_);
    and _3119_(_1331_, _1384_, packet_buffer_3[34]);
    and _3120_(_1332_, _1383_, packet_in[34]);
    or _3121_(_0328_, _1332_, _1331_);
    and _3122_(_1333_, _1384_, packet_buffer_3[35]);
    and _3123_(_1334_, _1383_, packet_in[35]);
    or _3124_(_0329_, _1334_, _1333_);
    and _3125_(_1335_, _1384_, packet_buffer_3[36]);
    and _3126_(_1336_, _1383_, packet_in[36]);
    or _3127_(_0330_, _1336_, _1335_);
    and _3128_(_1337_, _1384_, packet_buffer_3[37]);
    and _3129_(_1338_, _1383_, packet_in[37]);
    or _3130_(_0331_, _1338_, _1337_);
    and _3131_(_1339_, _1384_, packet_buffer_3[38]);
    and _3132_(_1340_, _1383_, packet_in[38]);
    or _3133_(_0332_, _1340_, _1339_);
    and _3134_(_1341_, _1384_, packet_buffer_3[39]);
    and _3135_(_1342_, _1383_, packet_in[39]);
    or _3136_(_0333_, _1342_, _1341_);
    and _3137_(_1343_, _1384_, packet_buffer_3[40]);
    and _3138_(_1344_, _1383_, packet_in[40]);
    or _3139_(_0334_, _1344_, _1343_);
    and _3140_(_1345_, _1384_, packet_buffer_3[41]);
    and _3141_(_1346_, _1383_, packet_in[41]);
    or _3142_(_0335_, _1346_, _1345_);
    and _3143_(_1347_, _1384_, packet_buffer_3[42]);
    and _3144_(_1348_, _1383_, packet_in[42]);
    or _3145_(_0336_, _1348_, _1347_);
    and _3146_(_1349_, _1384_, packet_buffer_3[43]);
    and _3147_(_1350_, _1383_, packet_in[43]);
    or _3148_(_0337_, _1350_, _1349_);
    and _3149_(_1351_, _1384_, packet_buffer_3[44]);
    and _3150_(_1352_, _1383_, packet_in[44]);
    or _3151_(_0338_, _1352_, _1351_);
    and _3152_(_1353_, _1384_, packet_buffer_3[45]);
    and _3153_(_1354_, _1383_, packet_in[45]);
    or _3154_(_0339_, _1354_, _1353_);
    and _3155_(_1355_, _1384_, packet_buffer_3[46]);
    and _3156_(_1356_, _1383_, packet_in[46]);
    or _3157_(_0340_, _1356_, _1355_);
    and _3158_(_1357_, _1384_, packet_buffer_3[47]);
    and _3159_(_1358_, _1383_, packet_in[47]);
    or _3160_(_0341_, _1358_, _1357_);
    and _3161_(_1359_, _1384_, packet_buffer_3[48]);
    and _3162_(_1360_, _1383_, packet_in[48]);
    or _3163_(_0342_, _1360_, _1359_);
    and _3164_(_1361_, _1384_, packet_buffer_3[49]);
    and _3165_(_1362_, _1383_, packet_in[49]);
    or _3166_(_0343_, _1362_, _1361_);
    and _3167_(_1363_, _1384_, packet_buffer_3[50]);
    and _3168_(_1364_, _1383_, packet_in[50]);
    or _3169_(_0344_, _1364_, _1363_);
    and _3170_(_1365_, _1384_, packet_buffer_3[51]);
    and _3171_(_1366_, _1383_, packet_in[51]);
    or _3172_(_0345_, _1366_, _1365_);
    xor _3173_(_0025_, _1410_, buffer_head[0]);
    xor _3174_(_1367_, buffer_head[1], buffer_head[0]);
    and _3175_(_1368_, _1367_, _1410_);
    nor _3176_(_1369_, _1410_, _1475_);
    or _3177_(_0026_, _1369_, _1368_);
    xor _3178_(_0027_, _1380_, buffer_tail[0]);
    xor _3179_(_1370_, buffer_tail[1], buffer_tail[0]);
    and _3180_(_1371_, _1370_, _1380_);
    nor _3181_(_1372_, _1380_, _0866_);
    or _3182_(_0028_, _1372_, _1371_);
    not _3183_(_1373_, packet_valid);
    nor _3184_(_1374_, _1447_, _1373_);
    and _3185_(_1375_, _1374_, _1450_);
    and _3186_(_1376_, _1451_, route_error);
    or _3187_(_0165_, _1376_, _1375_);
    not _3188_(_0001_, rst);
    not _3189_(_0002_, rst);
    not _3190_(_0003_, rst);
    not _3191_(_0004_, rst);
    not _3192_(_0005_, rst);
    not _3193_(_0006_, rst);
    not _3194_(_0007_, rst);
    not _3195_(_0008_, rst);
    not _3196_(_0009_, rst);
    not _3197_(_0010_, rst);
    not _3198_(_0011_, rst);
    not _3199_(_0012_, rst);
    dff _3200_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0013_), .Q(packet_buffer_3[52]));
    dff _3201_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0014_), .Q(packet_buffer_3[53]));
    dff _3202_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0015_), .Q(packet_buffer_3[54]));
    dff _3203_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0016_), .Q(packet_buffer_3[55]));
    dff _3204_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0017_), .Q(packet_buffer_3[56]));
    dff _3205_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0018_), .Q(packet_buffer_3[57]));
    dff _3206_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0019_), .Q(packet_buffer_3[58]));
    dff _3207_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0020_), .Q(packet_buffer_3[59]));
    dff _3208_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0021_), .Q(packet_buffer_3[60]));
    dff _3209_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0022_), .Q(packet_buffer_3[61]));
    dff _3210_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0023_), .Q(packet_buffer_3[62]));
    dff _3211_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0024_), .Q(packet_buffer_3[63]));
    dff _3212_(.RN(_0000_), .SN(1'b1), .CK(clk), .D(_0025_), .Q(buffer_head[0]));
    dff _3213_(.RN(_0001_), .SN(1'b1), .CK(clk), .D(_0026_), .Q(buffer_head[1]));
    dff _3214_(.RN(_0002_), .SN(1'b1), .CK(clk), .D(_0027_), .Q(buffer_tail[0]));
    dff _3215_(.RN(_0003_), .SN(1'b1), .CK(clk), .D(_0028_), .Q(buffer_tail[1]));
    dff _3216_(.RN(_0004_), .SN(1'b1), .CK(clk), .D(_0029_), .Q(packet_count[0]));
    dff _3217_(.RN(_0005_), .SN(1'b1), .CK(clk), .D(_0030_), .Q(packet_count[1]));
    dff _3218_(.RN(_0006_), .SN(1'b1), .CK(clk), .D(_0031_), .Q(packet_count[2]));
    dff _3219_(.RN(_0007_), .SN(1'b1), .CK(clk), .D(_0032_), .Q(packet_count[3]));
    dff _3220_(.RN(_0008_), .SN(1'b1), .CK(clk), .D(_0033_), .Q(network_state[0]));
    dff _3221_(.RN(_0009_), .SN(1'b1), .CK(clk), .D(_0034_), .Q(network_state[1]));
    dff _3222_(.RN(_0010_), .SN(1'b1), .CK(clk), .D(_0035_), .Q(network_state[2]));
    dff _3223_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0036_), .Q(packet_out[0]));
    dff _3224_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0037_), .Q(packet_out[1]));
    dff _3225_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0038_), .Q(packet_out[2]));
    dff _3226_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0039_), .Q(packet_out[3]));
    dff _3227_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0040_), .Q(packet_out[4]));
    dff _3228_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0041_), .Q(packet_out[5]));
    dff _3229_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0042_), .Q(packet_out[6]));
    dff _3230_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0043_), .Q(packet_out[7]));
    dff _3231_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0044_), .Q(packet_out[8]));
    dff _3232_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0045_), .Q(packet_out[9]));
    dff _3233_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0046_), .Q(packet_out[10]));
    dff _3234_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0047_), .Q(packet_out[11]));
    dff _3235_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0048_), .Q(packet_out[12]));
    dff _3236_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0049_), .Q(packet_out[13]));
    dff _3237_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0050_), .Q(packet_out[14]));
    dff _3238_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0051_), .Q(packet_out[15]));
    dff _3239_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0052_), .Q(packet_out[16]));
    dff _3240_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0053_), .Q(packet_out[17]));
    dff _3241_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0054_), .Q(packet_out[18]));
    dff _3242_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0055_), .Q(packet_out[19]));
    dff _3243_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0056_), .Q(packet_out[20]));
    dff _3244_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0057_), .Q(packet_out[21]));
    dff _3245_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0058_), .Q(packet_out[22]));
    dff _3246_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0059_), .Q(packet_out[23]));
    dff _3247_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0060_), .Q(packet_out[24]));
    dff _3248_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0061_), .Q(packet_out[25]));
    dff _3249_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0062_), .Q(packet_out[26]));
    dff _3250_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0063_), .Q(packet_out[27]));
    dff _3251_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0064_), .Q(packet_out[28]));
    dff _3252_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0065_), .Q(packet_out[29]));
    dff _3253_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0066_), .Q(packet_out[30]));
    dff _3254_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0067_), .Q(packet_out[31]));
    dff _3255_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0068_), .Q(packet_out[32]));
    dff _3256_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0069_), .Q(packet_out[33]));
    dff _3257_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0070_), .Q(packet_out[34]));
    dff _3258_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0071_), .Q(packet_out[35]));
    dff _3259_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0072_), .Q(packet_out[36]));
    dff _3260_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0073_), .Q(packet_out[37]));
    dff _3261_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0074_), .Q(packet_out[38]));
    dff _3262_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0075_), .Q(packet_out[39]));
    dff _3263_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0076_), .Q(packet_out[40]));
    dff _3264_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0077_), .Q(packet_out[41]));
    dff _3265_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0078_), .Q(packet_out[42]));
    dff _3266_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0079_), .Q(packet_out[43]));
    dff _3267_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0080_), .Q(packet_out[44]));
    dff _3268_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0081_), .Q(packet_out[45]));
    dff _3269_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0082_), .Q(packet_out[46]));
    dff _3270_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0083_), .Q(packet_out[47]));
    dff _3271_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0084_), .Q(packet_out[48]));
    dff _3272_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0085_), .Q(packet_out[49]));
    dff _3273_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0086_), .Q(packet_out[50]));
    dff _3274_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0087_), .Q(packet_out[51]));
    dff _3275_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0088_), .Q(packet_out[52]));
    dff _3276_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0089_), .Q(packet_out[53]));
    dff _3277_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0090_), .Q(packet_out[54]));
    dff _3278_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0091_), .Q(packet_out[55]));
    dff _3279_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0092_), .Q(packet_out[56]));
    dff _3280_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0093_), .Q(packet_out[57]));
    dff _3281_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0094_), .Q(packet_out[58]));
    dff _3282_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0095_), .Q(packet_out[59]));
    dff _3283_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0096_), .Q(packet_out[60]));
    dff _3284_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0097_), .Q(packet_out[61]));
    dff _3285_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0098_), .Q(packet_out[62]));
    dff _3286_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0099_), .Q(packet_out[63]));
    dff _3287_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0100_), .Q(packet_buffer_1[0]));
    dff _3288_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0101_), .Q(packet_buffer_1[1]));
    dff _3289_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0102_), .Q(packet_buffer_1[2]));
    dff _3290_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0103_), .Q(packet_buffer_1[3]));
    dff _3291_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0104_), .Q(packet_buffer_1[4]));
    dff _3292_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0105_), .Q(packet_buffer_1[5]));
    dff _3293_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0106_), .Q(packet_buffer_1[6]));
    dff _3294_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0107_), .Q(packet_buffer_1[7]));
    dff _3295_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0108_), .Q(packet_buffer_1[8]));
    dff _3296_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0109_), .Q(packet_buffer_1[9]));
    dff _3297_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0110_), .Q(packet_buffer_1[10]));
    dff _3298_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0111_), .Q(packet_buffer_1[11]));
    dff _3299_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0112_), .Q(packet_buffer_1[12]));
    dff _3300_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0113_), .Q(packet_buffer_1[13]));
    dff _3301_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0114_), .Q(packet_buffer_1[14]));
    dff _3302_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0115_), .Q(packet_buffer_1[15]));
    dff _3303_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0116_), .Q(packet_buffer_1[16]));
    dff _3304_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0117_), .Q(packet_buffer_1[17]));
    dff _3305_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0118_), .Q(packet_buffer_1[18]));
    dff _3306_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0119_), .Q(packet_buffer_1[19]));
    dff _3307_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0120_), .Q(packet_buffer_1[20]));
    dff _3308_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0121_), .Q(packet_buffer_1[21]));
    dff _3309_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0122_), .Q(packet_buffer_1[22]));
    dff _3310_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0123_), .Q(packet_buffer_1[23]));
    dff _3311_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0124_), .Q(packet_buffer_1[24]));
    dff _3312_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0125_), .Q(packet_buffer_1[25]));
    dff _3313_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0126_), .Q(packet_buffer_1[26]));
    dff _3314_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0127_), .Q(packet_buffer_1[27]));
    dff _3315_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0128_), .Q(packet_buffer_1[28]));
    dff _3316_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0129_), .Q(packet_buffer_1[29]));
    dff _3317_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0130_), .Q(packet_buffer_1[30]));
    dff _3318_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0131_), .Q(packet_buffer_1[31]));
    dff _3319_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0132_), .Q(packet_buffer_1[32]));
    dff _3320_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0133_), .Q(packet_buffer_1[33]));
    dff _3321_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0134_), .Q(packet_buffer_1[34]));
    dff _3322_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0135_), .Q(packet_buffer_1[35]));
    dff _3323_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0136_), .Q(packet_buffer_1[36]));
    dff _3324_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0137_), .Q(packet_buffer_1[37]));
    dff _3325_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0138_), .Q(packet_buffer_1[38]));
    dff _3326_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0139_), .Q(packet_buffer_1[39]));
    dff _3327_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0140_), .Q(packet_buffer_1[40]));
    dff _3328_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0141_), .Q(packet_buffer_1[41]));
    dff _3329_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0142_), .Q(packet_buffer_1[42]));
    dff _3330_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0143_), .Q(packet_buffer_1[43]));
    dff _3331_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0144_), .Q(packet_buffer_1[44]));
    dff _3332_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0145_), .Q(packet_buffer_1[45]));
    dff _3333_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0146_), .Q(packet_buffer_1[46]));
    dff _3334_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0147_), .Q(packet_buffer_1[47]));
    dff _3335_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0148_), .Q(packet_buffer_1[48]));
    dff _3336_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0149_), .Q(packet_buffer_1[49]));
    dff _3337_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0150_), .Q(packet_buffer_1[50]));
    dff _3338_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0151_), .Q(packet_buffer_1[51]));
    dff _3339_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0152_), .Q(packet_buffer_1[52]));
    dff _3340_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0153_), .Q(packet_buffer_1[53]));
    dff _3341_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0154_), .Q(packet_buffer_1[54]));
    dff _3342_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0155_), .Q(packet_buffer_1[55]));
    dff _3343_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0156_), .Q(packet_buffer_1[56]));
    dff _3344_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0157_), .Q(packet_buffer_1[57]));
    dff _3345_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0158_), .Q(packet_buffer_1[58]));
    dff _3346_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0159_), .Q(packet_buffer_1[59]));
    dff _3347_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0160_), .Q(packet_buffer_1[60]));
    dff _3348_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0161_), .Q(packet_buffer_1[61]));
    dff _3349_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0162_), .Q(packet_buffer_1[62]));
    dff _3350_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0163_), .Q(packet_buffer_1[63]));
    dff _3351_(.RN(_0011_), .SN(1'b1), .CK(clk), .D(_0164_), .Q(packet_ready));
    dff _3352_(.RN(_0012_), .SN(1'b1), .CK(clk), .D(_0165_), .Q(route_error));
    dff _3353_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0166_), .Q(packet_buffer_0[0]));
    dff _3354_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0167_), .Q(packet_buffer_0[1]));
    dff _3355_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0168_), .Q(packet_buffer_0[2]));
    dff _3356_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0169_), .Q(packet_buffer_0[3]));
    dff _3357_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0170_), .Q(packet_buffer_0[4]));
    dff _3358_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0171_), .Q(packet_buffer_0[5]));
    dff _3359_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0172_), .Q(packet_buffer_0[6]));
    dff _3360_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0173_), .Q(packet_buffer_0[7]));
    dff _3361_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0174_), .Q(packet_buffer_0[8]));
    dff _3362_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0175_), .Q(packet_buffer_0[9]));
    dff _3363_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0176_), .Q(packet_buffer_0[10]));
    dff _3364_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0177_), .Q(packet_buffer_0[11]));
    dff _3365_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0178_), .Q(packet_buffer_0[12]));
    dff _3366_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0179_), .Q(packet_buffer_0[13]));
    dff _3367_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0180_), .Q(packet_buffer_0[14]));
    dff _3368_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0181_), .Q(packet_buffer_0[15]));
    dff _3369_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0182_), .Q(packet_buffer_0[16]));
    dff _3370_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0183_), .Q(packet_buffer_0[17]));
    dff _3371_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0184_), .Q(packet_buffer_0[18]));
    dff _3372_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0185_), .Q(packet_buffer_0[19]));
    dff _3373_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0186_), .Q(packet_buffer_0[20]));
    dff _3374_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0187_), .Q(packet_buffer_0[21]));
    dff _3375_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0188_), .Q(packet_buffer_0[22]));
    dff _3376_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0189_), .Q(packet_buffer_0[23]));
    dff _3377_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0190_), .Q(packet_buffer_0[24]));
    dff _3378_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0191_), .Q(packet_buffer_0[25]));
    dff _3379_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0192_), .Q(packet_buffer_0[26]));
    dff _3380_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0193_), .Q(packet_buffer_0[27]));
    dff _3381_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0194_), .Q(packet_buffer_0[28]));
    dff _3382_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0195_), .Q(packet_buffer_0[29]));
    dff _3383_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0196_), .Q(packet_buffer_0[30]));
    dff _3384_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0197_), .Q(packet_buffer_0[31]));
    dff _3385_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0198_), .Q(packet_buffer_0[32]));
    dff _3386_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0199_), .Q(packet_buffer_0[33]));
    dff _3387_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0200_), .Q(packet_buffer_0[34]));
    dff _3388_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0201_), .Q(packet_buffer_0[35]));
    dff _3389_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0202_), .Q(packet_buffer_0[36]));
    dff _3390_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0203_), .Q(packet_buffer_0[37]));
    dff _3391_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0204_), .Q(packet_buffer_0[38]));
    dff _3392_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0205_), .Q(packet_buffer_0[39]));
    dff _3393_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0206_), .Q(packet_buffer_0[40]));
    dff _3394_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0207_), .Q(packet_buffer_0[41]));
    dff _3395_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0208_), .Q(packet_buffer_0[42]));
    dff _3396_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0209_), .Q(packet_buffer_0[43]));
    dff _3397_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0210_), .Q(packet_buffer_0[44]));
    dff _3398_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0211_), .Q(packet_buffer_0[45]));
    dff _3399_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0212_), .Q(packet_buffer_0[46]));
    dff _3400_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0213_), .Q(packet_buffer_0[47]));
    dff _3401_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0214_), .Q(packet_buffer_0[48]));
    dff _3402_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0215_), .Q(packet_buffer_0[49]));
    dff _3403_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0216_), .Q(packet_buffer_0[50]));
    dff _3404_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0217_), .Q(packet_buffer_0[51]));
    dff _3405_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0218_), .Q(packet_buffer_0[52]));
    dff _3406_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0219_), .Q(packet_buffer_0[53]));
    dff _3407_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0220_), .Q(packet_buffer_0[54]));
    dff _3408_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0221_), .Q(packet_buffer_0[55]));
    dff _3409_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0222_), .Q(packet_buffer_0[56]));
    dff _3410_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0223_), .Q(packet_buffer_0[57]));
    dff _3411_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0224_), .Q(packet_buffer_0[58]));
    dff _3412_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0225_), .Q(packet_buffer_0[59]));
    dff _3413_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0226_), .Q(packet_buffer_0[60]));
    dff _3414_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0227_), .Q(packet_buffer_0[61]));
    dff _3415_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0228_), .Q(packet_buffer_0[62]));
    dff _3416_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0229_), .Q(packet_buffer_0[63]));
    dff _3417_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0230_), .Q(packet_buffer_2[0]));
    dff _3418_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0231_), .Q(packet_buffer_2[1]));
    dff _3419_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0232_), .Q(packet_buffer_2[2]));
    dff _3420_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0233_), .Q(packet_buffer_2[3]));
    dff _3421_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0234_), .Q(packet_buffer_2[4]));
    dff _3422_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0235_), .Q(packet_buffer_2[5]));
    dff _3423_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0236_), .Q(packet_buffer_2[6]));
    dff _3424_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0237_), .Q(packet_buffer_2[7]));
    dff _3425_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0238_), .Q(packet_buffer_2[8]));
    dff _3426_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0239_), .Q(packet_buffer_2[9]));
    dff _3427_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0240_), .Q(packet_buffer_2[10]));
    dff _3428_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0241_), .Q(packet_buffer_2[11]));
    dff _3429_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0242_), .Q(packet_buffer_2[12]));
    dff _3430_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0243_), .Q(packet_buffer_2[13]));
    dff _3431_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0244_), .Q(packet_buffer_2[14]));
    dff _3432_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0245_), .Q(packet_buffer_2[15]));
    dff _3433_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0246_), .Q(packet_buffer_2[16]));
    dff _3434_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0247_), .Q(packet_buffer_2[17]));
    dff _3435_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0248_), .Q(packet_buffer_2[18]));
    dff _3436_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0249_), .Q(packet_buffer_2[19]));
    dff _3437_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0250_), .Q(packet_buffer_2[20]));
    dff _3438_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0251_), .Q(packet_buffer_2[21]));
    dff _3439_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0252_), .Q(packet_buffer_2[22]));
    dff _3440_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0253_), .Q(packet_buffer_2[23]));
    dff _3441_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0254_), .Q(packet_buffer_2[24]));
    dff _3442_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0255_), .Q(packet_buffer_2[25]));
    dff _3443_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0256_), .Q(packet_buffer_2[26]));
    dff _3444_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0257_), .Q(packet_buffer_2[27]));
    dff _3445_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0258_), .Q(packet_buffer_2[28]));
    dff _3446_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0259_), .Q(packet_buffer_2[29]));
    dff _3447_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0260_), .Q(packet_buffer_2[30]));
    dff _3448_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0261_), .Q(packet_buffer_2[31]));
    dff _3449_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0262_), .Q(packet_buffer_2[32]));
    dff _3450_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0263_), .Q(packet_buffer_2[33]));
    dff _3451_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0264_), .Q(packet_buffer_2[34]));
    dff _3452_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0265_), .Q(packet_buffer_2[35]));
    dff _3453_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0266_), .Q(packet_buffer_2[36]));
    dff _3454_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0267_), .Q(packet_buffer_2[37]));
    dff _3455_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0268_), .Q(packet_buffer_2[38]));
    dff _3456_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0269_), .Q(packet_buffer_2[39]));
    dff _3457_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0270_), .Q(packet_buffer_2[40]));
    dff _3458_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0271_), .Q(packet_buffer_2[41]));
    dff _3459_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0272_), .Q(packet_buffer_2[42]));
    dff _3460_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0273_), .Q(packet_buffer_2[43]));
    dff _3461_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0274_), .Q(packet_buffer_2[44]));
    dff _3462_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0275_), .Q(packet_buffer_2[45]));
    dff _3463_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0276_), .Q(packet_buffer_2[46]));
    dff _3464_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0277_), .Q(packet_buffer_2[47]));
    dff _3465_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0278_), .Q(packet_buffer_2[48]));
    dff _3466_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0279_), .Q(packet_buffer_2[49]));
    dff _3467_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0280_), .Q(packet_buffer_2[50]));
    dff _3468_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0281_), .Q(packet_buffer_2[51]));
    dff _3469_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0282_), .Q(packet_buffer_2[52]));
    dff _3470_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0283_), .Q(packet_buffer_2[53]));
    dff _3471_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0284_), .Q(packet_buffer_2[54]));
    dff _3472_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0285_), .Q(packet_buffer_2[55]));
    dff _3473_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0286_), .Q(packet_buffer_2[56]));
    dff _3474_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0287_), .Q(packet_buffer_2[57]));
    dff _3475_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0288_), .Q(packet_buffer_2[58]));
    dff _3476_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0289_), .Q(packet_buffer_2[59]));
    dff _3477_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0290_), .Q(packet_buffer_2[60]));
    dff _3478_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0291_), .Q(packet_buffer_2[61]));
    dff _3479_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0292_), .Q(packet_buffer_2[62]));
    dff _3480_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0293_), .Q(packet_buffer_2[63]));
    dff _3481_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0294_), .Q(packet_buffer_3[0]));
    dff _3482_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0295_), .Q(packet_buffer_3[1]));
    dff _3483_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0296_), .Q(packet_buffer_3[2]));
    dff _3484_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0297_), .Q(packet_buffer_3[3]));
    dff _3485_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0298_), .Q(packet_buffer_3[4]));
    dff _3486_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0299_), .Q(packet_buffer_3[5]));
    dff _3487_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0300_), .Q(packet_buffer_3[6]));
    dff _3488_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0301_), .Q(packet_buffer_3[7]));
    dff _3489_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0302_), .Q(packet_buffer_3[8]));
    dff _3490_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0303_), .Q(packet_buffer_3[9]));
    dff _3491_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0304_), .Q(packet_buffer_3[10]));
    dff _3492_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0305_), .Q(packet_buffer_3[11]));
    dff _3493_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0306_), .Q(packet_buffer_3[12]));
    dff _3494_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0307_), .Q(packet_buffer_3[13]));
    dff _3495_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0308_), .Q(packet_buffer_3[14]));
    dff _3496_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0309_), .Q(packet_buffer_3[15]));
    dff _3497_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0310_), .Q(packet_buffer_3[16]));
    dff _3498_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0311_), .Q(packet_buffer_3[17]));
    dff _3499_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0312_), .Q(packet_buffer_3[18]));
    dff _3500_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0313_), .Q(packet_buffer_3[19]));
    dff _3501_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0314_), .Q(packet_buffer_3[20]));
    dff _3502_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0315_), .Q(packet_buffer_3[21]));
    dff _3503_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0316_), .Q(packet_buffer_3[22]));
    dff _3504_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0317_), .Q(packet_buffer_3[23]));
    dff _3505_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0318_), .Q(packet_buffer_3[24]));
    dff _3506_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0319_), .Q(packet_buffer_3[25]));
    dff _3507_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0320_), .Q(packet_buffer_3[26]));
    dff _3508_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0321_), .Q(packet_buffer_3[27]));
    dff _3509_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0322_), .Q(packet_buffer_3[28]));
    dff _3510_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0323_), .Q(packet_buffer_3[29]));
    dff _3511_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0324_), .Q(packet_buffer_3[30]));
    dff _3512_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0325_), .Q(packet_buffer_3[31]));
    dff _3513_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0326_), .Q(packet_buffer_3[32]));
    dff _3514_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0327_), .Q(packet_buffer_3[33]));
    dff _3515_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0328_), .Q(packet_buffer_3[34]));
    dff _3516_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0329_), .Q(packet_buffer_3[35]));
    dff _3517_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0330_), .Q(packet_buffer_3[36]));
    dff _3518_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0331_), .Q(packet_buffer_3[37]));
    dff _3519_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0332_), .Q(packet_buffer_3[38]));
    dff _3520_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0333_), .Q(packet_buffer_3[39]));
    dff _3521_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0334_), .Q(packet_buffer_3[40]));
    dff _3522_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0335_), .Q(packet_buffer_3[41]));
    dff _3523_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0336_), .Q(packet_buffer_3[42]));
    dff _3524_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0337_), .Q(packet_buffer_3[43]));
    dff _3525_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0338_), .Q(packet_buffer_3[44]));
    dff _3526_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0339_), .Q(packet_buffer_3[45]));
    dff _3527_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0340_), .Q(packet_buffer_3[46]));
    dff _3528_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0341_), .Q(packet_buffer_3[47]));
    dff _3529_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0342_), .Q(packet_buffer_3[48]));
    dff _3530_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0343_), .Q(packet_buffer_3[49]));
    dff _3531_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0344_), .Q(packet_buffer_3[50]));
    dff _3532_(.RN(1'b1), .SN(1'b1), .CK(clk), .D(_0345_), .Q(packet_buffer_3[51]));
endmodule