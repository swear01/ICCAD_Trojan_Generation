module trojan0_rsa0_host_0000(clk, rst, message, modulus, exponent, rsa_start, result, rsa_done);
  wire _00000_;
  wire _00001_;
  wire _00002_;
  wire _00003_;
  wire _00004_;
  wire _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire [15:0] accumulator;
  wire [15:0] base;
  input clk;
  wire clk;
  wire [3:0] exp_counter;
  input [3:0] exponent;
  wire [3:0] exponent;
  input [15:0] message;
  wire [15:0] message;
  input [15:0] modulus;
  wire [15:0] modulus;
  output [15:0] result;
  wire [15:0] result;
  wire rsa_active;
  output rsa_done;
  wire rsa_done;
  input rsa_start;
  wire rsa_start;
  input rst;
  wire rst;
    not _06078_(_00001_, rst);
    not _06079_(_01138_, base[0]);
    not _06080_(_01149_, rsa_active);
    and _06081_(_01160_, rsa_start, _01149_);
    nor _06082_(_01171_, _01160_, _01149_);
    and _06083_(_01182_, base[14], base[1]);
    and _06084_(_01193_, base[15], base[0]);
    xnor _06085_(_01204_, _01193_, _01182_);
    and _06086_(_01215_, base[13], base[2]);
    xor _06087_(_01226_, _01215_, _01204_);
    nand _06088_(_01237_, base[13], base[1]);
    and _06089_(_01248_, base[14], base[0]);
    not _06090_(_01259_, _01248_);
    or _06091_(_01270_, _01259_, _01237_);
    and _06092_(_01281_, base[12], base[2]);
    not _06093_(_01292_, _01281_);
    xor _06094_(_01303_, _01248_, _01237_);
    or _06095_(_01314_, _01303_, _01292_);
    and _06096_(_01325_, _01314_, _01270_);
    xnor _06097_(_01336_, _01325_, _01226_);
    and _06098_(_01347_, base[12], base[3]);
    and _06099_(_01358_, base[11], base[4]);
    xnor _06100_(_01369_, _01358_, _01347_);
    and _06101_(_01380_, base[10], base[5]);
    xor _06102_(_01391_, _01380_, _01369_);
    xnor _06103_(_01402_, _01391_, _01336_);
    xor _06104_(_01413_, _01303_, _01281_);
    and _06105_(_01424_, base[12], base[1]);
    and _06106_(_01435_, base[13], base[0]);
    and _06107_(_01446_, _01435_, _01424_);
    not _06108_(_01457_, _01446_);
    and _06109_(_01468_, base[11], base[2]);
    not _06110_(_01479_, _01468_);
    xnor _06111_(_01490_, _01435_, _01424_);
    or _06112_(_01501_, _01490_, _01479_);
    and _06113_(_01512_, _01501_, _01457_);
    or _06114_(_01523_, _01512_, _01413_);
    and _06115_(_01534_, base[11], base[3]);
    and _06116_(_01545_, base[10], base[4]);
    xnor _06117_(_01556_, _01545_, _01534_);
    and _06118_(_01567_, base[9], base[5]);
    xor _06119_(_01578_, _01567_, _01556_);
    xnor _06120_(_01589_, _01512_, _01413_);
    or _06121_(_01600_, _01589_, _01578_);
    and _06122_(_01611_, _01600_, _01523_);
    xnor _06123_(_01622_, _01611_, _01402_);
    nand _06124_(_01633_, _01545_, _01534_);
    not _06125_(_01644_, _01567_);
    or _06126_(_01655_, _01644_, _01556_);
    and _06127_(_01666_, _01655_, _01633_);
    nand _06128_(_01687_, base[9], base[6]);
    xor _06129_(_01698_, _01687_, _01666_);
    and _06130_(_01709_, base[8], base[6]);
    nand _06131_(_01720_, _01709_, base[7]);
    not _06132_(_01731_, base[7]);
    nand _06133_(_01742_, _01709_, _01731_);
    and _06134_(_01753_, _01742_, _01720_);
    xor _06135_(_01764_, _01753_, _01698_);
    xnor _06136_(_01775_, _01764_, _01622_);
    xnor _06137_(_01786_, _01589_, _01578_);
    xor _06138_(_01797_, _01490_, _01468_);
    and _06139_(_01808_, base[11], base[1]);
    and _06140_(_01819_, base[12], base[0]);
    nand _06141_(_01830_, _01819_, _01808_);
    and _06142_(_01841_, base[10], base[2]);
    not _06143_(_01852_, _01841_);
    xnor _06144_(_01863_, _01819_, _01808_);
    or _06145_(_01874_, _01863_, _01852_);
    and _06146_(_01885_, _01874_, _01830_);
    or _06147_(_01896_, _01885_, _01797_);
    and _06148_(_01907_, base[9], base[4]);
    and _06149_(_01918_, base[10], base[3]);
    xnor _06150_(_01929_, _01918_, _01907_);
    and _06151_(_01940_, base[8], base[5]);
    xor _06152_(_01951_, _01940_, _01929_);
    xnor _06153_(_01962_, _01885_, _01797_);
    or _06154_(_01973_, _01962_, _01951_);
    and _06155_(_01984_, _01973_, _01896_);
    or _06156_(_01995_, _01984_, _01786_);
    and _06157_(_02006_, _01918_, _01907_);
    not _06158_(_02017_, _01940_);
    nor _06159_(_02028_, _02017_, _01929_);
    nor _06160_(_02039_, _02028_, _02006_);
    xnor _06161_(_02050_, _01709_, base[7]);
    xor _06162_(_02061_, _02050_, _01709_);
    xnor _06163_(_02072_, _02061_, _02039_);
    and _06164_(_02083_, base[7], base[6]);
    xor _06165_(_02094_, _02083_, _02072_);
    xnor _06166_(_02104_, _01984_, _01786_);
    or _06167_(_02114_, _02104_, _02094_);
    and _06168_(_02125_, _02114_, _01995_);
    xnor _06169_(_02136_, _02125_, _01775_);
    or _06170_(_02147_, _02061_, _02039_);
    not _06171_(_02158_, _02083_);
    or _06172_(_02169_, _02158_, _02072_);
    and _06173_(_02180_, _02169_, _02147_);
    nand _06174_(_02191_, base[9], base[6]);
    xor _06175_(_02202_, _02191_, _01380_);
    xor _06176_(_02213_, _02202_, _01358_);
    nand _06177_(_02224_, _01567_, _01545_);
    not _06178_(_02235_, _01534_);
    xnor _06179_(_02246_, _01567_, _01545_);
    or _06180_(_02257_, _02246_, _02235_);
    and _06181_(_02268_, _02257_, _02224_);
    xor _06182_(_02279_, _02268_, _02213_);
    xnor _06183_(_02290_, _01347_, _01215_);
    xor _06184_(_02301_, _02290_, _01182_);
    xor _06185_(_02312_, _02301_, _02279_);
    xor _06186_(_02323_, _02312_, _02180_);
    xor _06187_(_02334_, _02246_, _01534_);
    nor _06188_(_02345_, _01929_, _01479_);
    nor _06189_(_02356_, _02345_, _02006_);
    or _06190_(_02367_, _02356_, _02334_);
    xor _06191_(_02378_, _01281_, _01237_);
    xor _06192_(_02389_, _02378_, _01248_);
    xnor _06193_(_02400_, _02356_, _02334_);
    or _06194_(_02411_, _02400_, _02389_);
    and _06195_(_02422_, _02411_, _02367_);
    xor _06196_(_02433_, _02422_, _02323_);
    xnor _06197_(_02444_, _02433_, _02136_);
    xnor _06198_(_02455_, _02104_, _02094_);
    xnor _06199_(_02466_, _01962_, _01951_);
    xor _06200_(_02477_, _01863_, _01841_);
    and _06201_(_02488_, base[10], base[1]);
    and _06202_(_02499_, base[11], base[0]);
    nand _06203_(_02510_, _02499_, _02488_);
    and _06204_(_02521_, base[9], base[2]);
    not _06205_(_02532_, _02521_);
    xnor _06206_(_02543_, _02499_, _02488_);
    or _06207_(_02554_, _02543_, _02532_);
    and _06208_(_02565_, _02554_, _02510_);
    or _06209_(_02576_, _02565_, _02477_);
    and _06210_(_02587_, base[9], base[3]);
    and _06211_(_02598_, base[8], base[4]);
    xnor _06212_(_02609_, _02598_, _02587_);
    and _06213_(_02620_, base[7], base[5]);
    xor _06214_(_02631_, _02620_, _02609_);
    xnor _06215_(_02642_, _02565_, _02477_);
    or _06216_(_02653_, _02642_, _02631_);
    and _06217_(_02664_, _02653_, _02576_);
    or _06218_(_02675_, _02664_, _02466_);
    and _06219_(_02686_, _02598_, _02587_);
    not _06220_(_02697_, _02620_);
    nor _06221_(_02708_, _02697_, _02609_);
    nor _06222_(_02719_, _02708_, _02686_);
    xor _06223_(_02730_, _02719_, _01940_);
    and _06224_(_02741_, _02620_, base[6]);
    not _06225_(_02752_, _02598_);
    xnor _06226_(_02763_, _02620_, base[6]);
    nor _06227_(_02774_, _02763_, _02752_);
    nor _06228_(_02785_, _02774_, _02741_);
    xnor _06229_(_02796_, _02785_, _02730_);
    xnor _06230_(_02807_, _02664_, _02466_);
    or _06231_(_02818_, _02807_, _02796_);
    and _06232_(_02829_, _02818_, _02675_);
    or _06233_(_02840_, _02829_, _02455_);
    nor _06234_(_02851_, _02719_, _02017_);
    nor _06235_(_02862_, _02785_, _02730_);
    nor _06236_(_02873_, _02862_, _02851_);
    xnor _06237_(_02884_, _02400_, _02389_);
    xnor _06238_(_02895_, _02884_, _02873_);
    xor _06239_(_02906_, _01929_, _01468_);
    and _06240_(_02917_, _02587_, _01841_);
    not _06241_(_02928_, _01808_);
    xnor _06242_(_02939_, _02587_, _01841_);
    nor _06243_(_02950_, _02939_, _02928_);
    nor _06244_(_02961_, _02950_, _02917_);
    nor _06245_(_02972_, _02961_, _02906_);
    xnor _06246_(_02983_, _02961_, _02906_);
    nor _06247_(_02994_, _02983_, _01490_);
    nor _06248_(_03005_, _02994_, _02972_);
    xnor _06249_(_03016_, _03005_, _02895_);
    xnor _06250_(_03027_, _02829_, _02455_);
    or _06251_(_03038_, _03027_, _03016_);
    and _06252_(_03049_, _03038_, _02840_);
    xnor _06253_(_03060_, _03049_, _02444_);
    nor _06254_(_03071_, _02884_, _02873_);
    nor _06255_(_03082_, _03005_, _02895_);
    or _06256_(_03093_, _03082_, _03071_);
    or _06257_(_03104_, _01292_, _01237_);
    or _06258_(_03115_, _02378_, _01259_);
    and _06259_(_03126_, _03115_, _03104_);
    xor _06260_(_03137_, _03126_, _03093_);
    xor _06261_(_03148_, _03137_, _01193_);
    xnor _06262_(_03159_, _03148_, _03060_);
    xnor _06263_(_03170_, _03027_, _03016_);
    xnor _06264_(_03181_, _02807_, _02796_);
    xnor _06265_(_03192_, _02642_, _02631_);
    xor _06266_(_03203_, _02543_, _02521_);
    and _06267_(_03214_, base[9], base[1]);
    and _06268_(_03225_, base[10], base[0]);
    and _06269_(_03236_, _03225_, _03214_);
    not _06270_(_03247_, _03236_);
    and _06271_(_03258_, base[8], base[2]);
    not _06272_(_03269_, _03258_);
    xnor _06273_(_03280_, _03225_, _03214_);
    or _06274_(_03291_, _03280_, _03269_);
    and _06275_(_03302_, _03291_, _03247_);
    or _06276_(_03313_, _03302_, _03203_);
    and _06277_(_03324_, base[8], base[3]);
    and _06278_(_03335_, base[7], base[4]);
    xnor _06279_(_03346_, _03335_, _03324_);
    and _06280_(_03357_, base[6], base[5]);
    xor _06281_(_03368_, _03357_, _03346_);
    xnor _06282_(_03379_, _03302_, _03203_);
    or _06283_(_03390_, _03379_, _03368_);
    and _06284_(_03401_, _03390_, _03313_);
    or _06285_(_03412_, _03401_, _03192_);
    xor _06286_(_03423_, _02763_, _02598_);
    xnor _06287_(_03434_, _03401_, _03192_);
    or _06288_(_03445_, _03434_, _03423_);
    and _06289_(_03456_, _03445_, _03412_);
    or _06290_(_03467_, _03456_, _03181_);
    and _06291_(_03478_, _03335_, _03324_);
    not _06292_(_03489_, _03357_);
    nor _06293_(_03500_, _03489_, _03346_);
    nor _06294_(_03511_, _03500_, _03478_);
    xor _06295_(_03522_, _02763_, _02598_);
    nor _06296_(_03533_, _03522_, _03511_);
    xnor _06297_(_03544_, _03522_, _03511_);
    and _06298_(_03555_, _03357_, _03335_);
    not _06299_(_03566_, _03324_);
    xnor _06300_(_03577_, _03357_, _03335_);
    nor _06301_(_03588_, _03577_, _03566_);
    nor _06302_(_03599_, _03588_, _03555_);
    nor _06303_(_03610_, _03599_, _03544_);
    nor _06304_(_03621_, _03610_, _03533_);
    xnor _06305_(_03632_, _02983_, _01490_);
    xnor _06306_(_03643_, _03632_, _03621_);
    xor _06307_(_03654_, _02939_, _01808_);
    and _06308_(_03665_, _02521_, _02488_);
    not _06309_(_03676_, _02499_);
    xnor _06310_(_03687_, _02521_, _02488_);
    nor _06311_(_03698_, _03687_, _03676_);
    nor _06312_(_03709_, _03698_, _03665_);
    nor _06313_(_03720_, _03709_, _03654_);
    not _06314_(_03731_, _01819_);
    xnor _06315_(_03742_, _03709_, _03654_);
    nor _06316_(_03753_, _03742_, _03731_);
    nor _06317_(_03764_, _03753_, _03720_);
    xnor _06318_(_03775_, _03764_, _03643_);
    xnor _06319_(_03786_, _03456_, _03181_);
    or _06320_(_03797_, _03786_, _03775_);
    and _06321_(_03808_, _03797_, _03467_);
    or _06322_(_03819_, _03808_, _03170_);
    nor _06323_(_03830_, _03632_, _03621_);
    nor _06324_(_03841_, _03764_, _03643_);
    nor _06325_(_03852_, _03841_, _03830_);
    xor _06326_(_03863_, _03852_, _01446_);
    xnor _06327_(_03874_, _03808_, _03170_);
    or _06328_(_03885_, _03874_, _03863_);
    and _06329_(_03896_, _03885_, _03819_);
    xnor _06330_(_03907_, _03896_, _03159_);
    nor _06331_(_03918_, _03852_, _01457_);
    xor _06332_(_03929_, _03918_, _03907_);
    xnor _06333_(_03940_, _03874_, _03863_);
    xnor _06334_(_03951_, _03786_, _03775_);
    xnor _06335_(_03962_, _03434_, _03423_);
    xnor _06336_(_03973_, _03379_, _03368_);
    xor _06337_(_03984_, _03280_, _03258_);
    nand _06338_(_03995_, base[8], base[1]);
    and _06339_(_04006_, base[9], base[0]);
    not _06340_(_04017_, _04006_);
    or _06341_(_04028_, _04017_, _03995_);
    and _06342_(_04039_, base[7], base[2]);
    not _06343_(_04050_, _04039_);
    xor _06344_(_04061_, _04006_, _03995_);
    or _06345_(_04072_, _04061_, _04050_);
    and _06346_(_04083_, _04072_, _04028_);
    nor _06347_(_04094_, _04083_, _03984_);
    not _06348_(_04105_, _04094_);
    and _06349_(_04116_, base[6], base[4]);
    and _06350_(_04127_, base[7], base[3]);
    xnor _06351_(_04138_, _04127_, _04116_);
    xor _06352_(_04149_, _04138_, base[5]);
    xnor _06353_(_04160_, _04083_, _03984_);
    or _06354_(_04171_, _04160_, _04149_);
    and _06355_(_04182_, _04171_, _04105_);
    nor _06356_(_04193_, _04182_, _03973_);
    and _06357_(_04204_, _04127_, _04116_);
    not _06358_(_04215_, base[5]);
    nor _06359_(_04226_, _04138_, _04215_);
    nor _06360_(_04237_, _04226_, _04204_);
    xor _06361_(_04248_, _03577_, _03324_);
    xnor _06362_(_04259_, _04248_, _04237_);
    nor _06363_(_04270_, _04138_, _03269_);
    nor _06364_(_04281_, _04270_, _04204_);
    xnor _06365_(_04292_, _04281_, _04259_);
    xnor _06366_(_04303_, _04182_, _03973_);
    nor _06367_(_04314_, _04303_, _04292_);
    nor _06368_(_04325_, _04314_, _04193_);
    nor _06369_(_04336_, _04325_, _03962_);
    nor _06370_(_04347_, _04248_, _04237_);
    nor _06371_(_04358_, _04281_, _04259_);
    nor _06372_(_04369_, _04358_, _04347_);
    xor _06373_(_04380_, _03742_, _01819_);
    not _06374_(_04391_, _04380_);
    xor _06375_(_04402_, _04391_, _04369_);
    xor _06376_(_04413_, _03687_, _02499_);
    nor _06377_(_04424_, _04413_, _03247_);
    xor _06378_(_04435_, _04424_, _04402_);
    xnor _06379_(_04446_, _04325_, _03962_);
    nor _06380_(_04457_, _04446_, _04435_);
    nor _06381_(_04468_, _04457_, _04336_);
    nor _06382_(_04479_, _04468_, _03951_);
    nor _06383_(_04490_, _04380_, _04369_);
    not _06384_(_04501_, _04424_);
    nor _06385_(_04512_, _04501_, _04402_);
    nor _06386_(_04523_, _04512_, _04490_);
    xnor _06387_(_04534_, _04468_, _03951_);
    nor _06388_(_04545_, _04534_, _04523_);
    nor _06389_(_04556_, _04545_, _04479_);
    nor _06390_(_04567_, _04556_, _03940_);
    xor _06391_(_04578_, _04567_, _03929_);
    xnor _06392_(_04589_, _04556_, _03940_);
    not _06393_(_04600_, _04589_);
    xnor _06394_(_04611_, _04534_, _04523_);
    xnor _06395_(_04622_, _04446_, _04435_);
    xor _06396_(_04633_, _04303_, _04292_);
    not _06397_(_04644_, _04633_);
    xor _06398_(_04655_, _04160_, _04149_);
    not _06399_(_04666_, _04655_);
    xor _06400_(_04677_, _04061_, _04050_);
    not _06401_(_04688_, _04677_);
    nand _06402_(_04699_, base[7], base[1]);
    and _06403_(_04710_, base[8], base[0]);
    not _06404_(_04721_, _04710_);
    or _06405_(_04732_, _04721_, _04699_);
    and _06406_(_04743_, base[6], base[2]);
    not _06407_(_04754_, _04743_);
    xor _06408_(_04765_, _04710_, _04699_);
    or _06409_(_04776_, _04765_, _04754_);
    and _06410_(_04787_, _04776_, _04732_);
    or _06411_(_04798_, _04787_, _04688_);
    nand _06412_(_04819_, base[6], base[3]);
    xor _06413_(_04830_, _04787_, _04677_);
    or _06414_(_04841_, _04830_, _04819_);
    and _06415_(_04852_, _04841_, _04798_);
    or _06416_(_04863_, _04852_, _04666_);
    and _06417_(_04874_, base[6], base[3]);
    nand _06418_(_04885_, base[5], base[4]);
    xor _06419_(_04896_, _04138_, _03258_);
    xnor _06420_(_04907_, _04896_, _04885_);
    and _06421_(_04918_, _04874_, _04039_);
    xnor _06422_(_04929_, _04874_, _04039_);
    nor _06423_(_04940_, _04929_, _03995_);
    nor _06424_(_04951_, _04940_, _04918_);
    xnor _06425_(_04962_, _04951_, _04907_);
    xor _06426_(_04973_, _04852_, _04655_);
    or _06427_(_04984_, _04973_, _04962_);
    and _06428_(_04995_, _04984_, _04863_);
    nor _06429_(_05006_, _04995_, _04644_);
    not _06430_(_05017_, _05006_);
    nor _06431_(_05028_, _04896_, _04885_);
    nor _06432_(_05039_, _04951_, _04907_);
    nor _06433_(_05050_, _05039_, _05028_);
    xor _06434_(_05061_, _04413_, _03236_);
    xnor _06435_(_05072_, _05061_, _05050_);
    xor _06436_(_05083_, _04995_, _04633_);
    or _06437_(_05094_, _05083_, _05072_);
    and _06438_(_05105_, _05094_, _05017_);
    nor _06439_(_05116_, _05105_, _04622_);
    not _06440_(_05127_, _05116_);
    nor _06441_(_05138_, _05061_, _05050_);
    not _06442_(_05149_, _05138_);
    xnor _06443_(_05159_, _05105_, _04622_);
    or _06444_(_05169_, _05159_, _05149_);
    and _06445_(_05180_, _05169_, _05127_);
    nor _06446_(_05190_, _05180_, _04611_);
    nand _06447_(_05200_, _05190_, _04600_);
    xor _06448_(_05211_, _05190_, _04589_);
    xnor _06449_(_05221_, _05180_, _04611_);
    not _06450_(_05231_, _05221_);
    xor _06451_(_05242_, _05159_, _05138_);
    xor _06452_(_05252_, _05083_, _05072_);
    not _06453_(_05262_, _05252_);
    xnor _06454_(_05273_, _04973_, _04962_);
    xnor _06455_(_05283_, _04830_, _04819_);
    xor _06456_(_05293_, _04765_, _04743_);
    nand _06457_(_05304_, base[6], base[1]);
    not _06458_(_05314_, _05304_);
    and _06459_(_05324_, base[7], base[0]);
    nand _06460_(_05335_, _05324_, _05314_);
    and _06461_(_05345_, base[5], base[2]);
    not _06462_(_05355_, _05345_);
    xor _06463_(_05366_, _05324_, _05304_);
    or _06464_(_05376_, _05366_, _05355_);
    and _06465_(_05386_, _05376_, _05335_);
    or _06466_(_05397_, _05386_, _05293_);
    and _06467_(_05407_, base[5], base[3]);
    not _06468_(_05417_, base[4]);
    xor _06469_(_05428_, _05407_, _05417_);
    xor _06470_(_05438_, _05428_, _05407_);
    xnor _06471_(_05448_, _05386_, _05293_);
    or _06472_(_05459_, _05448_, _05438_);
    and _06473_(_05469_, _05459_, _05397_);
    or _06474_(_05480_, _05469_, _05283_);
    and _06475_(_05490_, _05407_, base[4]);
    and _06476_(_05500_, _05407_, _05417_);
    nor _06477_(_05511_, _05500_, _05490_);
    xnor _06478_(_05521_, _04929_, _03995_);
    xnor _06479_(_05532_, _05521_, _05511_);
    nor _06480_(_05542_, _04754_, _04699_);
    xor _06481_(_05552_, _04743_, _04699_);
    nor _06482_(_05563_, _05552_, _04721_);
    nor _06483_(_05573_, _05563_, _05542_);
    xnor _06484_(_05584_, _05573_, _05532_);
    xnor _06485_(_05594_, _05469_, _05283_);
    or _06486_(_05604_, _05594_, _05584_);
    and _06487_(_05615_, _05604_, _05480_);
    or _06488_(_05625_, _05615_, _05273_);
    nor _06489_(_05635_, _05521_, _05511_);
    nor _06490_(_05645_, _05573_, _05532_);
    nor _06491_(_05655_, _05645_, _05635_);
    xnor _06492_(_05664_, _05655_, _03280_);
    xnor _06493_(_05671_, _05615_, _05273_);
    or _06494_(_05679_, _05671_, _05664_);
    and _06495_(_05687_, _05679_, _05625_);
    nor _06496_(_05694_, _05687_, _05262_);
    nor _06497_(_05700_, _05655_, _03280_);
    not _06498_(_05701_, _05700_);
    xor _06499_(_05702_, _05687_, _05252_);
    nor _06500_(_05703_, _05702_, _05701_);
    nor _06501_(_05704_, _05703_, _05694_);
    nor _06502_(_05705_, _05704_, _05242_);
    nand _06503_(_05706_, _05705_, _05231_);
    xor _06504_(_05707_, _05705_, _05221_);
    xnor _06505_(_05708_, _05704_, _05242_);
    xor _06506_(_05709_, _05702_, _05701_);
    not _06507_(_05710_, _05709_);
    xnor _06508_(_05711_, _05671_, _05664_);
    xnor _06509_(_05712_, _05594_, _05584_);
    xnor _06510_(_05713_, _05448_, _05438_);
    xor _06511_(_05714_, _05366_, _05345_);
    nand _06512_(_05715_, base[5], base[1]);
    and _06513_(_05716_, base[6], base[0]);
    not _06514_(_05717_, _05716_);
    or _06515_(_05718_, _05717_, _05715_);
    and _06516_(_05719_, base[4], base[2]);
    not _06517_(_05720_, _05719_);
    xor _06518_(_05721_, _05716_, _05715_);
    or _06519_(_05722_, _05721_, _05720_);
    and _06520_(_05723_, _05722_, _05718_);
    or _06521_(_05724_, _05723_, _05714_);
    xnor _06522_(_05725_, _05723_, _05714_);
    or _06523_(_05726_, _05725_, _05355_);
    and _06524_(_05727_, _05726_, _05724_);
    or _06525_(_05728_, _05727_, _05713_);
    and _06526_(_05729_, base[4], base[3]);
    xor _06527_(_05730_, _05552_, _04710_);
    xor _06528_(_05731_, _05730_, _05729_);
    xnor _06529_(_05732_, _05731_, _05335_);
    xnor _06530_(_05733_, _05727_, _05713_);
    or _06531_(_05734_, _05733_, _05732_);
    and _06532_(_05735_, _05734_, _05728_);
    or _06533_(_05736_, _05735_, _05712_);
    not _06534_(_05737_, _05729_);
    nor _06535_(_05738_, _05730_, _05737_);
    nor _06536_(_05739_, _05731_, _05335_);
    nor _06537_(_05740_, _05739_, _05738_);
    xor _06538_(_05741_, _05740_, _04006_);
    xnor _06539_(_05742_, _05735_, _05712_);
    or _06540_(_05743_, _05742_, _05741_);
    and _06541_(_05744_, _05743_, _05736_);
    or _06542_(_05745_, _05744_, _05711_);
    nor _06543_(_05746_, _05740_, _04017_);
    not _06544_(_05747_, _05746_);
    xnor _06545_(_05748_, _05744_, _05711_);
    or _06546_(_05749_, _05748_, _05747_);
    and _06547_(_05750_, _05749_, _05745_);
    or _06548_(_05751_, _05750_, _05710_);
    or _06549_(_05752_, _05751_, _05708_);
    or _06550_(_05753_, _05752_, _05707_);
    and _06551_(_05754_, _05753_, _05706_);
    xnor _06552_(_05755_, _05751_, _05708_);
    or _06553_(_05756_, _05755_, _05707_);
    xor _06554_(_05757_, _05750_, _05709_);
    xor _06555_(_05758_, _05748_, _05747_);
    xnor _06556_(_05759_, _05742_, _05741_);
    xnor _06557_(_05760_, _05733_, _05732_);
    xor _06558_(_05761_, _05725_, _05345_);
    xor _06559_(_05762_, _05721_, _05719_);
    nand _06560_(_05763_, base[4], base[1]);
    and _06561_(_05764_, base[5], base[0]);
    not _06562_(_05765_, _05764_);
    or _06563_(_05766_, _05765_, _05763_);
    and _06564_(_05767_, base[3], base[2]);
    not _06565_(_05768_, _05767_);
    xor _06566_(_05769_, _05764_, _05763_);
    or _06567_(_05770_, _05769_, _05768_);
    and _06568_(_05771_, _05770_, _05766_);
    or _06569_(_05772_, _05771_, _05762_);
    not _06570_(_05773_, base[3]);
    xor _06571_(_05774_, _05719_, _05773_);
    xnor _06572_(_05775_, _05774_, _05715_);
    xnor _06573_(_05776_, _05771_, _05762_);
    or _06574_(_05777_, _05776_, _05775_);
    and _06575_(_05778_, _05777_, _05772_);
    or _06576_(_05779_, _05778_, _05761_);
    and _06577_(_05780_, _05719_, base[3]);
    nor _06578_(_05781_, _05774_, _05715_);
    nor _06579_(_05782_, _05781_, _05780_);
    xnor _06580_(_05783_, _05782_, _05366_);
    xnor _06581_(_05784_, _05778_, _05761_);
    or _06582_(_05785_, _05784_, _05783_);
    and _06583_(_05786_, _05785_, _05779_);
    or _06584_(_05787_, _05786_, _05760_);
    nor _06585_(_05788_, _05782_, _05366_);
    not _06586_(_05789_, _05788_);
    xnor _06587_(_05790_, _05786_, _05760_);
    or _06588_(_05791_, _05790_, _05789_);
    and _06589_(_05792_, _05791_, _05787_);
    nor _06590_(_05793_, _05792_, _05759_);
    nand _06591_(_05794_, _05793_, _05758_);
    or _06592_(_05795_, _05794_, _05757_);
    xnor _06593_(_05796_, _05794_, _05757_);
    xnor _06594_(_05797_, _05793_, _05758_);
    xor _06595_(_05798_, _05792_, _05759_);
    xor _06596_(_05799_, _05790_, _05788_);
    xnor _06597_(_05800_, _05784_, _05783_);
    xnor _06598_(_05801_, _05776_, _05775_);
    xor _06599_(_05802_, _05769_, _05767_);
    nand _06600_(_05803_, base[3], base[1]);
    nand _06601_(_05804_, base[4], base[0]);
    or _06602_(_05805_, _05804_, _05803_);
    not _06603_(_05806_, base[2]);
    xnor _06604_(_05807_, _05804_, _05803_);
    or _06605_(_05808_, _05807_, _05806_);
    and _06606_(_05809_, _05808_, _05805_);
    or _06607_(_05810_, _05809_, _05802_);
    xor _06608_(_05811_, _05767_, _05763_);
    xor _06609_(_05812_, _05811_, _05764_);
    xnor _06610_(_05813_, _05809_, _05802_);
    or _06611_(_05814_, _05813_, _05812_);
    and _06612_(_05815_, _05814_, _05810_);
    or _06613_(_05816_, _05815_, _05801_);
    nor _06614_(_05817_, _05768_, _05763_);
    nor _06615_(_05818_, _05811_, _05765_);
    nor _06616_(_05819_, _05818_, _05817_);
    xor _06617_(_05820_, _05819_, _05716_);
    xnor _06618_(_05821_, _05815_, _05801_);
    or _06619_(_05822_, _05821_, _05820_);
    and _06620_(_05823_, _05822_, _05816_);
    or _06621_(_05824_, _05823_, _05800_);
    nor _06622_(_05825_, _05819_, _05717_);
    not _06623_(_05826_, _05825_);
    xnor _06624_(_05827_, _05823_, _05800_);
    or _06625_(_05828_, _05827_, _05826_);
    and _06626_(_05829_, _05828_, _05824_);
    nor _06627_(_05830_, _05829_, _05799_);
    nand _06628_(_05831_, _05830_, _05798_);
    or _06629_(_05832_, _05831_, _05797_);
    or _06630_(_05833_, _05832_, _05796_);
    and _06631_(_05834_, _05833_, _05795_);
    xnor _06632_(_05835_, _05831_, _05797_);
    or _06633_(_05836_, _05835_, _05796_);
    xnor _06634_(_05837_, _05830_, _05798_);
    xor _06635_(_05838_, _05829_, _05799_);
    xor _06636_(_05839_, _05827_, _05826_);
    xnor _06637_(_05840_, _05821_, _05820_);
    xnor _06638_(_05841_, _05813_, _05812_);
    xor _06639_(_05842_, _05807_, base[2]);
    and _06640_(_05843_, base[3], base[0]);
    nand _06641_(_05844_, base[2], base[1]);
    nor _06642_(_05845_, _05844_, _05842_);
    and _06643_(_05846_, base[2], base[1]);
    xor _06644_(_05847_, _05846_, _05842_);
    nor _06645_(_05848_, _05847_, _05807_);
    nor _06646_(_05849_, _05848_, _05845_);
    nor _06647_(_05850_, _05849_, _05841_);
    xnor _06648_(_05851_, _05849_, _05841_);
    nor _06649_(_05852_, _05851_, _05805_);
    nor _06650_(_05853_, _05852_, _05850_);
    nor _06651_(_05854_, _05853_, _05840_);
    and _06652_(_05855_, _05854_, _05839_);
    nand _06653_(_05856_, _05855_, _05838_);
    or _06654_(_05857_, _05856_, _05837_);
    xnor _06655_(_05858_, _05856_, _05837_);
    xnor _06656_(_05859_, _05855_, _05838_);
    xor _06657_(_05860_, _05854_, _05839_);
    xnor _06658_(_05861_, _05853_, _05840_);
    not _06659_(_05862_, _05861_);
    xnor _06660_(_05863_, _05851_, _05805_);
    or _06661_(_05864_, _05806_, base[1]);
    not _06662_(_05865_, base[1]);
    nand _06663_(_05866_, base[2], base[0]);
    or _06664_(_05867_, _05866_, _05865_);
    or _06665_(_05868_, _05866_, base[1]);
    and _06666_(_05869_, _05868_, _05867_);
    nand _06667_(_05870_, base[3], base[0]);
    nor _06668_(_05871_, _05870_, _05864_);
    not _06669_(_05872_, _05871_);
    nor _06670_(_05873_, _05872_, _05863_);
    nand _06671_(_05874_, _05873_, _05862_);
    not _06672_(_05875_, _05874_);
    nand _06673_(_05876_, _05875_, _05860_);
    or _06674_(_05877_, _05876_, _05859_);
    or _06675_(_05878_, _05877_, _05858_);
    and _06676_(_05879_, _05878_, _05857_);
    or _06677_(_05880_, _05879_, _05836_);
    and _06678_(_05881_, _05880_, _05834_);
    xnor _06679_(_05882_, _05876_, _05859_);
    or _06680_(_05883_, _05882_, _05858_);
    or _06681_(_05884_, _05883_, _05836_);
    xor _06682_(_05885_, _05874_, _05860_);
    not _06683_(_05886_, _05885_);
    xor _06684_(_05887_, _05873_, _05861_);
    xnor _06685_(_05888_, _05871_, _05863_);
    xor _06686_(_05889_, _05870_, _05864_);
    and _06687_(_05890_, base[3], base[0]);
    xor _06688_(_05891_, _05869_, _05890_);
    xor _06689_(_05892_, _05891_, _05843_);
    nand _06690_(_05893_, base[1], base[0]);
    nor _06691_(_05894_, _05893_, _05892_);
    and _06692_(_05895_, _05894_, _05889_);
    and _06693_(_05896_, _05895_, _05888_);
    not _06694_(_05897_, _05896_);
    nor _06695_(_05898_, _05897_, _05887_);
    and _06696_(_05899_, _05898_, _05886_);
    not _06697_(_05900_, _05899_);
    or _06698_(_05901_, _05900_, _05884_);
    and _06699_(_05902_, _05901_, _05881_);
    or _06700_(_05903_, _05902_, _05756_);
    and _06701_(_05904_, _05903_, _05754_);
    or _06702_(_05905_, _05904_, _05211_);
    and _06703_(_05906_, _05905_, _05200_);
    xnor _06704_(_05907_, _05906_, _04578_);
    or _06705_(_05908_, _05900_, _05883_);
    and _06706_(_05909_, _05908_, _05879_);
    or _06707_(_05910_, _05909_, _05835_);
    and _06708_(_05911_, _05910_, _05832_);
    xnor _06709_(_05912_, _05911_, _05796_);
    xnor _06710_(_05913_, _05909_, _05835_);
    and _06711_(_05914_, _05913_, _05912_);
    or _06712_(_05915_, _05900_, _05882_);
    and _06713_(_05916_, _05915_, _05877_);
    xnor _06714_(_05917_, _05916_, _05858_);
    xor _06715_(_05918_, _05899_, _05882_);
    and _06716_(_05919_, _05918_, _05917_);
    and _06717_(_05920_, _05919_, _05914_);
    not _06718_(_05921_, _05920_);
    or _06719_(_05922_, _05902_, _05755_);
    and _06720_(_05923_, _05922_, _05752_);
    xnor _06721_(_05924_, _05923_, _05707_);
    xnor _06722_(_05925_, _05902_, _05755_);
    nand _06723_(_05926_, _05925_, _05924_);
    not _06724_(_05927_, modulus[0]);
    xor _06725_(_05928_, _05907_, _05927_);
    xnor _06726_(_05929_, _05904_, _05211_);
    not _06727_(_05930_, _05929_);
    or _06728_(_05931_, _05930_, _05928_);
    or _06729_(_05932_, _05931_, _05926_);
    or _06730_(_05933_, _05932_, _05921_);
    xor _06731_(_05934_, _05898_, _05885_);
    xor _06732_(_05935_, _05896_, _05887_);
    and _06733_(_05936_, _05935_, _05934_);
    xor _06734_(_05937_, _05895_, _05888_);
    xnor _06735_(_05938_, _05894_, _05889_);
    not _06736_(_05939_, _05938_);
    nor _06737_(_05940_, _05939_, _05937_);
    and _06738_(_05941_, _05940_, _05936_);
    nor _06739_(_05942_, base[1], base[0]);
    and _06740_(_05943_, _05942_, _05941_);
    not _06741_(_05944_, _05943_);
    nor _06742_(_05945_, _05944_, _05933_);
    nor _06743_(_05946_, modulus[8], modulus[7]);
    nor _06744_(_05947_, modulus[6], modulus[5]);
    and _06745_(_05948_, _05947_, _05946_);
    nor _06746_(_05949_, modulus[2], modulus[1]);
    nor _06747_(_05950_, modulus[4], modulus[3]);
    and _06748_(_05951_, _05950_, _05949_);
    and _06749_(_05952_, _05951_, _05948_);
    nor _06750_(_05953_, modulus[12], modulus[11]);
    nor _06751_(_05954_, modulus[10], modulus[9]);
    and _06752_(_05955_, _05954_, _05953_);
    not _06753_(_05956_, modulus[15]);
    nor _06754_(_05957_, modulus[14], modulus[13]);
    and _06755_(_05958_, _05957_, _05956_);
    and _06756_(_05959_, _05958_, _05955_);
    and _06757_(_05960_, _05959_, _05952_);
    nand _06758_(_05961_, _05960_, _05945_);
    or _06759_(_05962_, _05907_, modulus[0]);
    or _06760_(_05963_, _05929_, _05928_);
    and _06761_(_05964_, _05963_, _05962_);
    and _06762_(_05965_, _05925_, _05924_);
    or _06763_(_05966_, _05965_, _05931_);
    and _06764_(_05967_, _05966_, _05964_);
    and _06765_(_05968_, _05913_, _05912_);
    not _06766_(_05969_, _05968_);
    and _06767_(_05970_, _05918_, _05917_);
    not _06768_(_05971_, _05970_);
    and _06769_(_05972_, _05971_, _05914_);
    nor _06770_(_05973_, _05972_, _05969_);
    or _06771_(_05974_, _05973_, _05932_);
    and _06772_(_05975_, _05974_, _05967_);
    and _06773_(_05976_, _05935_, _05934_);
    or _06774_(_05977_, _05939_, _05937_);
    nand _06775_(_05978_, _05977_, _05936_);
    and _06776_(_05979_, _05978_, _05976_);
    xnor _06777_(_05980_, _05893_, _05892_);
    or _06778_(_05981_, _05865_, base[0]);
    nand _06779_(_05982_, _05940_, _05936_);
    and _06780_(_05983_, _05982_, _05979_);
    or _06781_(_05984_, _05983_, _05933_);
    nand _06782_(_05985_, _05984_, _05975_);
    and _06783_(_05986_, _05985_, _05952_);
    and _06784_(_05987_, _05986_, _05955_);
    and _06785_(_05988_, _05987_, _05957_);
    nand _06786_(_05989_, _05988_, _05956_);
    nand _06787_(_05990_, _05989_, _05961_);
    or _06788_(_05991_, _05990_, _05907_);
    and _06789_(_05992_, _05989_, _05961_);
    not _06790_(_05993_, _05983_);
    nand _06791_(_05994_, _05993_, _05920_);
    and _06792_(_05995_, _05994_, _05973_);
    or _06793_(_05996_, _05995_, _05926_);
    and _06794_(_05997_, _05996_, _05965_);
    nand _06795_(_05998_, _05997_, _05929_);
    xor _06796_(_05999_, _05998_, _05928_);
    or _06797_(_06000_, _05999_, _05992_);
    and _06798_(_06001_, _06000_, _05991_);
    or _06799_(_06002_, _05990_, _05912_);
    nand _06800_(_06003_, _05993_, _05919_);
    and _06801_(_06004_, _06003_, _05970_);
    and _06802_(_06005_, _06004_, _05913_);
    xor _06803_(_06006_, _06005_, _05912_);
    or _06804_(_06007_, _06006_, _05992_);
    nand _06805_(_06008_, _06007_, _06002_);
    or _06806_(_06009_, _05990_, _05913_);
    xor _06807_(_06010_, _06004_, _05913_);
    or _06808_(_06011_, _06010_, _05992_);
    nand _06809_(_06012_, _06011_, _06009_);
    or _06810_(_06013_, _06012_, _06008_);
    or _06811_(_06014_, _05990_, _05917_);
    and _06812_(_06015_, _05983_, _05918_);
    xor _06813_(_06016_, _06015_, _05917_);
    or _06814_(_06017_, _06016_, _05992_);
    and _06815_(_06018_, _06017_, _06014_);
    or _06816_(_06019_, _05990_, _05918_);
    xor _06817_(_06020_, _05983_, _05918_);
    or _06818_(_06021_, _06020_, _05992_);
    and _06819_(_06022_, _06021_, _06019_);
    nand _06820_(_06023_, _06022_, _06018_);
    or _06821_(_06024_, _06023_, _06013_);
    or _06822_(_06025_, _05990_, _05924_);
    and _06823_(_06026_, _05995_, _05925_);
    xor _06824_(_06027_, _06026_, _05924_);
    or _06825_(_06028_, _06027_, _05992_);
    and _06826_(_06029_, _06028_, _06025_);
    or _06827_(_06030_, _05990_, _05925_);
    xor _06828_(_06031_, _05995_, _05925_);
    or _06829_(_06032_, _06031_, _05992_);
    and _06830_(_06033_, _06032_, _06030_);
    nand _06831_(_06034_, _06033_, _06029_);
    not _06832_(_06035_, modulus[1]);
    xor _06833_(_06036_, _06001_, _06035_);
    or _06834_(_06037_, _05990_, _05929_);
    xor _06835_(_06038_, _05997_, _05929_);
    or _06836_(_06039_, _06038_, _05992_);
    and _06837_(_06040_, _06039_, _06037_);
    xor _06838_(_06041_, _06040_, _05927_);
    or _06839_(_06042_, _06041_, _06036_);
    or _06840_(_06043_, _06042_, _06034_);
    or _06841_(_06044_, _06043_, _06024_);
    not _06842_(_06045_, _05942_);
    or _06843_(_06046_, _05990_, _05934_);
    nor _06844_(_06047_, _05939_, _05937_);
    nor _06845_(_06048_, _06047_, _05977_);
    and _06846_(_06049_, _06048_, _05935_);
    xor _06847_(_06050_, _06049_, _05934_);
    or _06848_(_06051_, _06050_, _05992_);
    nand _06849_(_06052_, _06051_, _06046_);
    or _06850_(_06053_, _05990_, _05935_);
    xor _06851_(_06054_, _06048_, _05935_);
    or _06852_(_06055_, _06054_, _05992_);
    nand _06853_(_06056_, _06055_, _06053_);
    or _06854_(_06057_, _06056_, _06052_);
    nor _06855_(_06058_, _05939_, _05937_);
    not _06856_(_06059_, _06058_);
    or _06857_(_06060_, _06059_, _06057_);
    nor _06858_(_06061_, _06060_, _06045_);
    not _06859_(_06062_, _06061_);
    nor _06860_(_06063_, _06062_, _06044_);
    nor _06861_(_06064_, modulus[3], modulus[2]);
    nor _06862_(_06065_, modulus[5], modulus[4]);
    and _06863_(_06066_, _06065_, _06064_);
    nor _06864_(_06067_, modulus[9], modulus[8]);
    nor _06865_(_06068_, modulus[7], modulus[6]);
    and _06866_(_06069_, _06068_, _06067_);
    and _06867_(_06070_, _06069_, _06066_);
    nor _06868_(_06071_, modulus[14], modulus[15]);
    nor _06869_(_06072_, modulus[10], modulus[11]);
    nor _06870_(_06073_, modulus[13], modulus[12]);
    and _06871_(_06074_, _06073_, _06072_);
    and _06872_(_06075_, _06074_, _06071_);
    and _06873_(_06076_, _06075_, _06070_);
    nand _06874_(_06077_, _06076_, _06063_);
    or _06875_(_00108_, _06001_, modulus[1]);
    or _06876_(_00109_, _06040_, modulus[0]);
    or _06877_(_00110_, _00109_, _06036_);
    and _06878_(_00111_, _00110_, _00108_);
    and _06879_(_00112_, _06033_, _06029_);
    or _06880_(_00113_, _00112_, _06042_);
    and _06881_(_00114_, _00113_, _00111_);
    nor _06882_(_00115_, _06012_, _06008_);
    and _06883_(_00116_, _06022_, _06018_);
    or _06884_(_00117_, _00116_, _06013_);
    and _06885_(_00118_, _00117_, _00115_);
    or _06886_(_00119_, _00118_, _06043_);
    and _06887_(_00120_, _00119_, _00114_);
    nor _06888_(_00121_, _06056_, _06052_);
    nor _06889_(_00122_, _05939_, _05937_);
    or _06890_(_00123_, _00122_, _06057_);
    and _06891_(_00124_, _00123_, _00121_);
    and _06892_(_00125_, _05981_, _05980_);
    not _06893_(_00126_, _00125_);
    and _06894_(_00127_, _05981_, _05980_);
    and _06895_(_00128_, _00127_, _00126_);
    or _06896_(_00129_, _06060_, _00128_);
    and _06897_(_00130_, _00129_, _00124_);
    or _06898_(_00131_, _00130_, _06044_);
    nand _06899_(_00132_, _00131_, _00120_);
    and _06900_(_00133_, _00132_, _06070_);
    and _06901_(_00134_, _00133_, _06074_);
    nand _06902_(_00135_, _00134_, _06071_);
    nand _06903_(_00136_, _00135_, _06077_);
    or _06904_(_00137_, _00136_, _06001_);
    not _06905_(_00138_, _00136_);
    or _06906_(_00139_, _00130_, _06024_);
    and _06907_(_00140_, _00139_, _00118_);
    or _06908_(_00141_, _00140_, _06034_);
    and _06909_(_00142_, _00141_, _00112_);
    or _06910_(_00143_, _00142_, _06041_);
    nand _06911_(_00144_, _00143_, _00109_);
    xor _06912_(_00145_, _00144_, _06036_);
    or _06913_(_00146_, _00145_, _00138_);
    and _06914_(_00147_, _00146_, _00137_);
    nand _06915_(_00148_, _00138_, _06008_);
    not _06916_(_00149_, _06012_);
    or _06917_(_00150_, _00130_, _06023_);
    and _06918_(_00151_, _00150_, _00116_);
    and _06919_(_00152_, _00151_, _00149_);
    xor _06920_(_00153_, _00152_, _06008_);
    nand _06921_(_00154_, _00153_, _00136_);
    nand _06922_(_00155_, _00154_, _00148_);
    or _06923_(_00156_, _00136_, _00149_);
    xor _06924_(_00157_, _00151_, _00149_);
    or _06925_(_00158_, _00157_, _00138_);
    nand _06926_(_00159_, _00158_, _00156_);
    or _06927_(_00160_, _00159_, _00155_);
    or _06928_(_00161_, _00136_, _06018_);
    and _06929_(_00162_, _00130_, _06022_);
    xor _06930_(_00163_, _00162_, _06018_);
    or _06931_(_00164_, _00163_, _00138_);
    and _06932_(_00165_, _00164_, _00161_);
    or _06933_(_00166_, _00136_, _06022_);
    xor _06934_(_00167_, _00130_, _06022_);
    or _06935_(_00168_, _00167_, _00138_);
    and _06936_(_00169_, _00168_, _00166_);
    nand _06937_(_00170_, _00169_, _00165_);
    or _06938_(_00171_, _00170_, _00160_);
    or _06939_(_00172_, _00136_, _06029_);
    nand _06940_(_00173_, _00140_, _06033_);
    xor _06941_(_00174_, _00173_, _06029_);
    nand _06942_(_00175_, _00174_, _00136_);
    and _06943_(_00176_, _00175_, _00172_);
    xor _06944_(_00177_, _00176_, modulus[0]);
    or _06945_(_00178_, _00136_, _06033_);
    xor _06946_(_00179_, _00140_, _06033_);
    or _06947_(_00180_, _00179_, _00138_);
    and _06948_(_00181_, _00180_, _00178_);
    nand _06949_(_00182_, _00181_, _00177_);
    not _06950_(_00183_, modulus[2]);
    xor _06951_(_00184_, _00147_, _00183_);
    or _06952_(_00185_, _00136_, _06040_);
    xor _06953_(_00186_, _00142_, _06041_);
    nand _06954_(_00187_, _00186_, _00136_);
    and _06955_(_00188_, _00187_, _00185_);
    xor _06956_(_00189_, _00188_, _06035_);
    or _06957_(_00190_, _00189_, _00184_);
    or _06958_(_00191_, _00190_, _00182_);
    or _06959_(_00192_, _00191_, _00171_);
    not _06960_(_00193_, _06052_);
    or _06961_(_00194_, _00136_, _00193_);
    not _06962_(_00195_, _06056_);
    or _06963_(_00196_, _05939_, _05937_);
    and _06964_(_00197_, _00196_, _00122_);
    and _06965_(_00198_, _00197_, _00195_);
    xor _06966_(_00199_, _00198_, _00193_);
    or _06967_(_00200_, _00199_, _00138_);
    nand _06968_(_00201_, _00200_, _00194_);
    or _06969_(_00202_, _00136_, _00195_);
    xnor _06970_(_00203_, _00197_, _06056_);
    or _06971_(_00204_, _00203_, _00138_);
    nand _06972_(_00205_, _00204_, _00202_);
    or _06973_(_00206_, _00205_, _00201_);
    nand _06974_(_00207_, _05992_, _05937_);
    xnor _06975_(_00208_, _05895_, _05888_);
    or _06976_(_00209_, _00208_, _05992_);
    and _06977_(_00210_, _00209_, _00207_);
    or _06978_(_00211_, _00136_, _00210_);
    xnor _06979_(_00212_, _05894_, _05889_);
    and _06980_(_00213_, _00212_, _00128_);
    xor _06981_(_00214_, _00213_, _00210_);
    or _06982_(_00215_, _00214_, _00138_);
    and _06983_(_00216_, _00215_, _00211_);
    or _06984_(_00217_, _00136_, _00212_);
    xor _06985_(_00218_, _05894_, _05889_);
    nand _06986_(_00219_, _00218_, _00136_);
    and _06987_(_00220_, _00219_, _00217_);
    nand _06988_(_00221_, _00220_, _00216_);
    or _06989_(_00222_, _00221_, _00206_);
    nor _06990_(_00223_, _00222_, _06045_);
    not _06991_(_00224_, _00223_);
    nor _06992_(_00225_, _00224_, _00192_);
    and _06993_(_00226_, _05954_, _05946_);
    and _06994_(_00227_, _05950_, _05947_);
    and _06995_(_00228_, _00227_, _00226_);
    and _06996_(_00229_, _05957_, _05953_);
    and _06997_(_00230_, _00229_, _05956_);
    and _06998_(_00231_, _00230_, _00228_);
    nand _06999_(_00232_, _00231_, _00225_);
    or _07000_(_00233_, _00147_, modulus[2]);
    or _07001_(_00234_, _00188_, modulus[1]);
    or _07002_(_00235_, _00234_, _00184_);
    and _07003_(_00236_, _00235_, _00233_);
    or _07004_(_00237_, _00176_, modulus[0]);
    xor _07005_(_00238_, _00176_, _05927_);
    or _07006_(_00239_, _00181_, _00238_);
    and _07007_(_00240_, _00239_, _00237_);
    or _07008_(_00241_, _00240_, _00190_);
    and _07009_(_00242_, _00241_, _00236_);
    nor _07010_(_00243_, _00159_, _00155_);
    and _07011_(_00244_, _00169_, _00165_);
    or _07012_(_00245_, _00244_, _00160_);
    and _07013_(_00246_, _00245_, _00243_);
    or _07014_(_00247_, _00246_, _00191_);
    and _07015_(_00248_, _00247_, _00242_);
    nor _07016_(_00249_, _00205_, _00201_);
    and _07017_(_00250_, _00220_, _00216_);
    or _07018_(_00251_, _00250_, _00206_);
    and _07019_(_00252_, _00251_, _00249_);
    or _07020_(_00253_, _00222_, _00128_);
    and _07021_(_00254_, _00253_, _00252_);
    or _07022_(_00255_, _00254_, _00192_);
    nand _07023_(_00256_, _00255_, _00248_);
    and _07024_(_00257_, _00256_, _00228_);
    and _07025_(_00258_, _00257_, _00229_);
    nand _07026_(_00259_, _00258_, _05956_);
    nand _07027_(_00260_, _00259_, _00232_);
    or _07028_(_00261_, _00260_, _00147_);
    and _07029_(_00262_, _00259_, _00232_);
    or _07030_(_00263_, _00254_, _00171_);
    and _07031_(_00264_, _00263_, _00246_);
    or _07032_(_00265_, _00264_, _00182_);
    and _07033_(_00266_, _00265_, _00240_);
    or _07034_(_00267_, _00266_, _00189_);
    nand _07035_(_00268_, _00267_, _00234_);
    xor _07036_(_00269_, _00268_, _00184_);
    or _07037_(_00270_, _00269_, _00262_);
    and _07038_(_00271_, _00270_, _00261_);
    not _07039_(_00272_, _00155_);
    or _07040_(_00273_, _00260_, _00272_);
    not _07041_(_00274_, _00159_);
    or _07042_(_00275_, _00254_, _00170_);
    and _07043_(_00276_, _00275_, _00244_);
    and _07044_(_00277_, _00276_, _00274_);
    xor _07045_(_00278_, _00277_, _00272_);
    or _07046_(_00279_, _00278_, _00262_);
    and _07047_(_00280_, _00279_, _00273_);
    or _07048_(_00281_, _00260_, _00274_);
    xor _07049_(_00282_, _00276_, _00274_);
    or _07050_(_00283_, _00282_, _00262_);
    and _07051_(_00284_, _00283_, _00281_);
    nand _07052_(_00285_, _00284_, _00280_);
    or _07053_(_00286_, _00260_, _00165_);
    and _07054_(_00287_, _00254_, _00169_);
    xor _07055_(_00288_, _00287_, _00165_);
    or _07056_(_00289_, _00288_, _00262_);
    and _07057_(_00290_, _00289_, _00286_);
    or _07058_(_00291_, _00260_, _00169_);
    xor _07059_(_00292_, _00254_, _00169_);
    or _07060_(_00293_, _00292_, _00262_);
    and _07061_(_00294_, _00293_, _00291_);
    nand _07062_(_00295_, _00294_, _00290_);
    or _07063_(_00296_, _00295_, _00285_);
    or _07064_(_00297_, _00260_, _00176_);
    and _07065_(_00298_, _00264_, _00181_);
    xnor _07066_(_00299_, _00298_, _00238_);
    or _07067_(_00300_, _00299_, _00262_);
    and _07068_(_00301_, _00300_, _00297_);
    xor _07069_(_00302_, _00301_, _06035_);
    or _07070_(_00303_, _00260_, _00181_);
    xor _07071_(_00304_, _00264_, _00181_);
    or _07072_(_00305_, _00304_, _00262_);
    and _07073_(_00306_, _00305_, _00303_);
    xor _07074_(_00307_, _00306_, _05927_);
    or _07075_(_00308_, _00307_, _00302_);
    not _07076_(_00309_, modulus[3]);
    xor _07077_(_00310_, _00271_, _00309_);
    or _07078_(_00311_, _00260_, _00188_);
    xnor _07079_(_00312_, _00266_, _00189_);
    or _07080_(_00313_, _00312_, _00262_);
    and _07081_(_00314_, _00313_, _00311_);
    xor _07082_(_00315_, _00314_, _00183_);
    or _07083_(_00316_, _00315_, _00310_);
    or _07084_(_00317_, _00316_, _00308_);
    nor _07085_(_00318_, _00317_, _00296_);
    not _07086_(_00319_, _00201_);
    or _07087_(_00320_, _00260_, _00319_);
    not _07088_(_00321_, _00205_);
    or _07089_(_00322_, _00221_, _00128_);
    and _07090_(_00323_, _00322_, _00250_);
    and _07091_(_00324_, _00323_, _00321_);
    xor _07092_(_00325_, _00324_, _00319_);
    or _07093_(_00326_, _00325_, _00262_);
    nand _07094_(_00327_, _00326_, _00320_);
    or _07095_(_00328_, _00260_, _00321_);
    xor _07096_(_00329_, _00323_, _00321_);
    or _07097_(_00330_, _00329_, _00262_);
    nand _07098_(_00331_, _00330_, _00328_);
    or _07099_(_00332_, _00331_, _00327_);
    or _07100_(_00333_, _00260_, _00216_);
    and _07101_(_00334_, _00220_, _00128_);
    xor _07102_(_00335_, _00334_, _00216_);
    or _07103_(_00336_, _00335_, _00262_);
    and _07104_(_00337_, _00336_, _00333_);
    or _07105_(_00338_, _00260_, _00220_);
    xor _07106_(_00339_, _00220_, _00128_);
    or _07107_(_00340_, _00339_, _00262_);
    and _07108_(_00341_, _00340_, _00338_);
    nand _07109_(_00342_, _00341_, _00337_);
    nor _07110_(_00343_, _00342_, _00332_);
    and _07111_(_00344_, _00343_, _05942_);
    and _07112_(_00345_, _00344_, _00318_);
    and _07113_(_00346_, _06073_, _06071_);
    and _07114_(_00347_, _06072_, _06067_);
    and _07115_(_00348_, _06068_, _06065_);
    and _07116_(_00349_, _00348_, _00347_);
    and _07117_(_00350_, _00349_, _00346_);
    nand _07118_(_00351_, _00350_, _00345_);
    or _07119_(_00352_, _00271_, modulus[3]);
    or _07120_(_00353_, _00314_, modulus[2]);
    or _07121_(_00354_, _00353_, _00310_);
    and _07122_(_00355_, _00354_, _00352_);
    or _07123_(_00356_, _00301_, modulus[1]);
    or _07124_(_00357_, _00306_, modulus[0]);
    or _07125_(_00358_, _00357_, _00302_);
    and _07126_(_00359_, _00358_, _00356_);
    or _07127_(_00360_, _00359_, _00316_);
    and _07128_(_00361_, _00360_, _00355_);
    and _07129_(_00362_, _00284_, _00280_);
    and _07130_(_00363_, _00294_, _00290_);
    or _07131_(_00364_, _00363_, _00285_);
    and _07132_(_00365_, _00364_, _00362_);
    or _07133_(_00366_, _00365_, _00317_);
    and _07134_(_00367_, _00366_, _00361_);
    nor _07135_(_00368_, _00331_, _00327_);
    and _07136_(_00369_, _00341_, _00337_);
    or _07137_(_00370_, _00369_, _00332_);
    and _07138_(_00371_, _00370_, _00368_);
    not _07139_(_00372_, _00128_);
    nand _07140_(_00373_, _00343_, _00372_);
    and _07141_(_00374_, _00373_, _00371_);
    not _07142_(_00375_, _00374_);
    nand _07143_(_00376_, _00375_, _00318_);
    nand _07144_(_00377_, _00376_, _00367_);
    and _07145_(_00378_, _00377_, _00349_);
    nand _07146_(_00379_, _00378_, _00346_);
    nand _07147_(_00380_, _00379_, _00351_);
    or _07148_(_00381_, _00380_, _00271_);
    or _07149_(_00382_, _00374_, _00296_);
    and _07150_(_00383_, _00382_, _00365_);
    or _07151_(_00384_, _00383_, _00308_);
    and _07152_(_00385_, _00384_, _00359_);
    or _07153_(_00386_, _00385_, _00315_);
    and _07154_(_00387_, _00386_, _00353_);
    xor _07155_(_00388_, _00387_, _00310_);
    nand _07156_(_00389_, _00388_, _00380_);
    and _07157_(_00390_, _00389_, _00381_);
    or _07158_(_00391_, _00380_, _00280_);
    or _07159_(_00392_, _00374_, _00295_);
    and _07160_(_00393_, _00392_, _00363_);
    nand _07161_(_00394_, _00393_, _00284_);
    xor _07162_(_00395_, _00394_, _00280_);
    nand _07163_(_00396_, _00395_, _00380_);
    and _07164_(_00397_, _00396_, _00391_);
    xor _07165_(_00398_, _00397_, _05927_);
    or _07166_(_00399_, _00380_, _00284_);
    not _07167_(_00400_, _00380_);
    xor _07168_(_00401_, _00393_, _00284_);
    or _07169_(_00402_, _00401_, _00400_);
    nand _07170_(_00403_, _00402_, _00399_);
    or _07171_(_00404_, _00403_, _00398_);
    or _07172_(_00405_, _00380_, _00290_);
    and _07173_(_00406_, _00374_, _00294_);
    xor _07174_(_00407_, _00406_, _00290_);
    or _07175_(_00408_, _00407_, _00400_);
    and _07176_(_00409_, _00408_, _00405_);
    or _07177_(_00410_, _00380_, _00294_);
    xor _07178_(_00411_, _00374_, _00294_);
    or _07179_(_00412_, _00411_, _00400_);
    and _07180_(_00413_, _00412_, _00410_);
    nand _07181_(_00414_, _00413_, _00409_);
    or _07182_(_00415_, _00414_, _00404_);
    or _07183_(_00416_, _00380_, _00301_);
    or _07184_(_00417_, _00383_, _00307_);
    and _07185_(_00418_, _00417_, _00357_);
    xor _07186_(_00419_, _00418_, _00302_);
    nand _07187_(_00420_, _00419_, _00380_);
    and _07188_(_00421_, _00420_, _00416_);
    xor _07189_(_00422_, _00421_, _00183_);
    or _07190_(_00423_, _00380_, _00306_);
    xor _07191_(_00424_, _00383_, _00307_);
    nand _07192_(_00425_, _00424_, _00380_);
    and _07193_(_00426_, _00425_, _00423_);
    xor _07194_(_00427_, _00426_, _06035_);
    or _07195_(_00428_, _00427_, _00422_);
    not _07196_(_00429_, modulus[4]);
    xor _07197_(_00430_, _00390_, _00429_);
    or _07198_(_00431_, _00380_, _00314_);
    xor _07199_(_00432_, _00385_, _00315_);
    nand _07200_(_00433_, _00432_, _00380_);
    and _07201_(_00434_, _00433_, _00431_);
    xor _07202_(_00435_, _00434_, _00309_);
    or _07203_(_00436_, _00435_, _00430_);
    or _07204_(_00437_, _00436_, _00428_);
    nor _07205_(_00438_, _00437_, _00415_);
    not _07206_(_00439_, _00327_);
    or _07207_(_00440_, _00380_, _00439_);
    not _07208_(_00441_, _00331_);
    or _07209_(_00442_, _00342_, _00128_);
    and _07210_(_00443_, _00442_, _00369_);
    and _07211_(_00444_, _00443_, _00441_);
    xor _07212_(_00445_, _00444_, _00439_);
    or _07213_(_00446_, _00445_, _00400_);
    nand _07214_(_00447_, _00446_, _00440_);
    or _07215_(_00448_, _00380_, _00441_);
    xor _07216_(_00449_, _00443_, _00441_);
    or _07217_(_00450_, _00449_, _00400_);
    nand _07218_(_00451_, _00450_, _00448_);
    or _07219_(_00452_, _00451_, _00447_);
    or _07220_(_00453_, _00380_, _00337_);
    and _07221_(_00454_, _00341_, _00128_);
    xor _07222_(_00455_, _00454_, _00337_);
    or _07223_(_00456_, _00455_, _00400_);
    and _07224_(_00457_, _00456_, _00453_);
    or _07225_(_00458_, _00380_, _00341_);
    xor _07226_(_00459_, _00341_, _00128_);
    or _07227_(_00460_, _00459_, _00400_);
    and _07228_(_00461_, _00460_, _00458_);
    nand _07229_(_00462_, _00461_, _00457_);
    nor _07230_(_00463_, _00462_, _00452_);
    and _07231_(_00464_, _00463_, _05942_);
    and _07232_(_00465_, _00464_, _00438_);
    and _07233_(_00466_, _05955_, _05948_);
    and _07234_(_00467_, _00466_, _05958_);
    nand _07235_(_00468_, _00467_, _00465_);
    or _07236_(_00469_, _00390_, modulus[4]);
    or _07237_(_00470_, _00434_, modulus[3]);
    or _07238_(_00471_, _00470_, _00430_);
    and _07239_(_00472_, _00471_, _00469_);
    or _07240_(_00473_, _00421_, modulus[2]);
    or _07241_(_00474_, _00426_, modulus[1]);
    or _07242_(_00475_, _00474_, _00422_);
    and _07243_(_00476_, _00475_, _00473_);
    or _07244_(_00477_, _00476_, _00436_);
    and _07245_(_00478_, _00477_, _00472_);
    or _07246_(_00479_, _00397_, modulus[0]);
    and _07247_(_00480_, _00402_, _00399_);
    or _07248_(_00481_, _00480_, _00398_);
    and _07249_(_00482_, _00481_, _00479_);
    and _07250_(_00483_, _00413_, _00409_);
    or _07251_(_00484_, _00483_, _00404_);
    and _07252_(_00485_, _00484_, _00482_);
    or _07253_(_00486_, _00485_, _00437_);
    and _07254_(_00487_, _00486_, _00478_);
    nor _07255_(_00488_, _00451_, _00447_);
    and _07256_(_00489_, _00461_, _00457_);
    or _07257_(_00490_, _00489_, _00452_);
    and _07258_(_00491_, _00490_, _00488_);
    nand _07259_(_00492_, _00463_, _00372_);
    nand _07260_(_00493_, _00492_, _00491_);
    nand _07261_(_00494_, _00493_, _00438_);
    nand _07262_(_00495_, _00494_, _00487_);
    and _07263_(_00496_, _00495_, _00466_);
    and _07264_(_00497_, _00496_, _05957_);
    nand _07265_(_00498_, _00497_, _05956_);
    nand _07266_(_00499_, _00498_, _00468_);
    or _07267_(_00500_, _00499_, _00390_);
    and _07268_(_00501_, _00492_, _00491_);
    or _07269_(_00502_, _00501_, _00415_);
    and _07270_(_00503_, _00502_, _00485_);
    or _07271_(_00504_, _00503_, _00428_);
    and _07272_(_00505_, _00504_, _00476_);
    or _07273_(_00506_, _00505_, _00435_);
    and _07274_(_00507_, _00506_, _00470_);
    xor _07275_(_00508_, _00507_, _00430_);
    nand _07276_(_00509_, _00508_, _00499_);
    and _07277_(_00510_, _00509_, _00500_);
    or _07278_(_00511_, _00499_, _00397_);
    and _07279_(_00512_, _00498_, _00468_);
    or _07280_(_00513_, _00501_, _00414_);
    and _07281_(_00514_, _00513_, _00483_);
    and _07282_(_00515_, _00514_, _00480_);
    xnor _07283_(_00516_, _00515_, _00398_);
    or _07284_(_00517_, _00516_, _00512_);
    and _07285_(_00518_, _00517_, _00511_);
    xor _07286_(_00519_, _00518_, _06035_);
    or _07287_(_00520_, _00499_, _00480_);
    xor _07288_(_00521_, _00514_, _00480_);
    or _07289_(_00522_, _00521_, _00512_);
    and _07290_(_00523_, _00522_, _00520_);
    xor _07291_(_00524_, _00523_, _05927_);
    or _07292_(_00525_, _00524_, _00519_);
    or _07293_(_00526_, _00499_, _00409_);
    and _07294_(_00527_, _00501_, _00413_);
    xor _07295_(_00528_, _00527_, _00409_);
    or _07296_(_00529_, _00528_, _00512_);
    and _07297_(_00530_, _00529_, _00526_);
    or _07298_(_00531_, _00499_, _00413_);
    xor _07299_(_00532_, _00501_, _00413_);
    or _07300_(_00533_, _00532_, _00512_);
    and _07301_(_00534_, _00533_, _00531_);
    nand _07302_(_00535_, _00534_, _00530_);
    or _07303_(_00536_, _00535_, _00525_);
    or _07304_(_00537_, _00499_, _00421_);
    or _07305_(_00538_, _00503_, _00427_);
    and _07306_(_00539_, _00538_, _00474_);
    xor _07307_(_00540_, _00539_, _00422_);
    nand _07308_(_00541_, _00540_, _00499_);
    and _07309_(_00542_, _00541_, _00537_);
    xor _07310_(_00543_, _00542_, _00309_);
    or _07311_(_00544_, _00499_, _00426_);
    xnor _07312_(_00545_, _00503_, _00427_);
    or _07313_(_00546_, _00545_, _00512_);
    and _07314_(_00547_, _00546_, _00544_);
    xor _07315_(_00548_, _00547_, _00183_);
    or _07316_(_00549_, _00548_, _00543_);
    not _07317_(_00550_, modulus[5]);
    xor _07318_(_00551_, _00510_, _00550_);
    or _07319_(_00552_, _00499_, _00434_);
    xor _07320_(_00553_, _00505_, _00435_);
    nand _07321_(_00554_, _00553_, _00499_);
    and _07322_(_00555_, _00554_, _00552_);
    xor _07323_(_00556_, _00555_, _00429_);
    or _07324_(_00557_, _00556_, _00551_);
    or _07325_(_00558_, _00557_, _00549_);
    nor _07326_(_00559_, _00558_, _00536_);
    not _07327_(_00560_, _00447_);
    or _07328_(_00561_, _00499_, _00560_);
    not _07329_(_00562_, _00451_);
    or _07330_(_00563_, _00462_, _00128_);
    and _07331_(_00564_, _00563_, _00489_);
    and _07332_(_00565_, _00564_, _00562_);
    xor _07333_(_00566_, _00565_, _00560_);
    or _07334_(_00567_, _00566_, _00512_);
    and _07335_(_00568_, _00567_, _00561_);
    or _07336_(_00569_, _00499_, _00562_);
    xor _07337_(_00570_, _00564_, _00562_);
    or _07338_(_00571_, _00570_, _00512_);
    and _07339_(_00572_, _00571_, _00569_);
    nand _07340_(_00573_, _00572_, _00568_);
    or _07341_(_00574_, _00499_, _00457_);
    and _07342_(_00575_, _00461_, _00128_);
    xor _07343_(_00576_, _00575_, _00457_);
    or _07344_(_00577_, _00576_, _00512_);
    and _07345_(_00578_, _00577_, _00574_);
    or _07346_(_00579_, _00499_, _00461_);
    xor _07347_(_00580_, _00461_, _00128_);
    or _07348_(_00581_, _00580_, _00512_);
    and _07349_(_00582_, _00581_, _00579_);
    nand _07350_(_00583_, _00582_, _00578_);
    nor _07351_(_00584_, _00583_, _00573_);
    and _07352_(_00585_, _00584_, _05942_);
    and _07353_(_00586_, _00585_, _00559_);
    and _07354_(_00587_, _06074_, _06069_);
    and _07355_(_00588_, _00587_, _06071_);
    nand _07356_(_00589_, _00588_, _00586_);
    or _07357_(_00590_, _00510_, modulus[5]);
    or _07358_(_00591_, _00555_, modulus[4]);
    or _07359_(_00592_, _00591_, _00551_);
    and _07360_(_00593_, _00592_, _00590_);
    or _07361_(_00594_, _00542_, modulus[3]);
    or _07362_(_00595_, _00547_, modulus[2]);
    or _07363_(_00596_, _00595_, _00543_);
    and _07364_(_00597_, _00596_, _00594_);
    or _07365_(_00598_, _00597_, _00557_);
    and _07366_(_00599_, _00598_, _00593_);
    or _07367_(_00600_, _00518_, modulus[1]);
    or _07368_(_00601_, _00523_, modulus[0]);
    or _07369_(_00602_, _00601_, _00519_);
    and _07370_(_00603_, _00602_, _00600_);
    and _07371_(_00604_, _00534_, _00530_);
    or _07372_(_00605_, _00604_, _00525_);
    and _07373_(_00606_, _00605_, _00603_);
    or _07374_(_00607_, _00606_, _00558_);
    and _07375_(_00608_, _00607_, _00599_);
    and _07376_(_00609_, _00572_, _00568_);
    and _07377_(_00610_, _00582_, _00578_);
    or _07378_(_00611_, _00610_, _00573_);
    and _07379_(_00612_, _00611_, _00609_);
    nand _07380_(_00613_, _00584_, _00372_);
    and _07381_(_00614_, _00613_, _00612_);
    not _07382_(_00615_, _00614_);
    nand _07383_(_00616_, _00615_, _00559_);
    nand _07384_(_00617_, _00616_, _00608_);
    and _07385_(_00618_, _00617_, _00587_);
    nand _07386_(_00619_, _00618_, _06071_);
    nand _07387_(_00620_, _00619_, _00589_);
    or _07388_(_00621_, _00620_, _00510_);
    or _07389_(_00622_, _00614_, _00536_);
    and _07390_(_00623_, _00622_, _00606_);
    or _07391_(_00624_, _00623_, _00549_);
    and _07392_(_00625_, _00624_, _00597_);
    or _07393_(_00626_, _00625_, _00556_);
    and _07394_(_00627_, _00626_, _00591_);
    xor _07395_(_00628_, _00627_, _00551_);
    nand _07396_(_00629_, _00628_, _00620_);
    and _07397_(_00630_, _00629_, _00621_);
    or _07398_(_00631_, _00620_, _00518_);
    or _07399_(_00632_, _00614_, _00535_);
    and _07400_(_00633_, _00632_, _00604_);
    or _07401_(_00634_, _00633_, _00524_);
    and _07402_(_00635_, _00634_, _00601_);
    xor _07403_(_00636_, _00635_, _00519_);
    nand _07404_(_00637_, _00636_, _00620_);
    and _07405_(_00638_, _00637_, _00631_);
    xor _07406_(_00639_, _00638_, _00183_);
    or _07407_(_00640_, _00620_, _00523_);
    and _07408_(_00641_, _00619_, _00589_);
    xnor _07409_(_00642_, _00633_, _00524_);
    or _07410_(_00643_, _00642_, _00641_);
    and _07411_(_00644_, _00643_, _00640_);
    xor _07412_(_00645_, _00644_, _06035_);
    or _07413_(_00646_, _00645_, _00639_);
    or _07414_(_00647_, _00620_, _00530_);
    and _07415_(_00648_, _00614_, _00534_);
    xor _07416_(_00649_, _00648_, _00530_);
    or _07417_(_00650_, _00649_, _00641_);
    and _07418_(_00651_, _00650_, _00647_);
    xor _07419_(_00652_, _00651_, _05927_);
    or _07420_(_00653_, _00620_, _00534_);
    xor _07421_(_00654_, _00614_, _00534_);
    or _07422_(_00655_, _00654_, _00641_);
    and _07423_(_00656_, _00655_, _00653_);
    not _07424_(_00657_, _00656_);
    or _07425_(_00658_, _00657_, _00652_);
    or _07426_(_00659_, _00658_, _00646_);
    or _07427_(_00660_, _00620_, _00542_);
    or _07428_(_00661_, _00623_, _00548_);
    and _07429_(_00662_, _00661_, _00595_);
    xor _07430_(_00663_, _00662_, _00543_);
    nand _07431_(_00664_, _00663_, _00620_);
    and _07432_(_00665_, _00664_, _00660_);
    xor _07433_(_00666_, _00665_, _00429_);
    or _07434_(_00667_, _00620_, _00547_);
    xnor _07435_(_00668_, _00623_, _00548_);
    or _07436_(_00669_, _00668_, _00641_);
    and _07437_(_00670_, _00669_, _00667_);
    xor _07438_(_00671_, _00670_, _00309_);
    or _07439_(_00672_, _00671_, _00666_);
    not _07440_(_00673_, modulus[6]);
    xor _07441_(_00674_, _00630_, _00673_);
    or _07442_(_00675_, _00620_, _00555_);
    xor _07443_(_00676_, _00625_, _00556_);
    nand _07444_(_00677_, _00676_, _00620_);
    and _07445_(_00678_, _00677_, _00675_);
    xor _07446_(_00679_, _00678_, _00550_);
    or _07447_(_00680_, _00679_, _00674_);
    or _07448_(_00681_, _00680_, _00672_);
    nor _07449_(_00682_, _00681_, _00659_);
    or _07450_(_00683_, _00620_, _00568_);
    or _07451_(_00684_, _00583_, _00128_);
    and _07452_(_00685_, _00684_, _00610_);
    and _07453_(_00686_, _00685_, _00572_);
    xor _07454_(_00687_, _00686_, _00568_);
    or _07455_(_00688_, _00687_, _00641_);
    and _07456_(_00689_, _00688_, _00683_);
    or _07457_(_00690_, _00620_, _00572_);
    xor _07458_(_00691_, _00685_, _00572_);
    or _07459_(_00692_, _00691_, _00641_);
    and _07460_(_00693_, _00692_, _00690_);
    nand _07461_(_00694_, _00693_, _00689_);
    or _07462_(_00695_, _00620_, _00578_);
    and _07463_(_00696_, _00582_, _00128_);
    xor _07464_(_00697_, _00696_, _00578_);
    or _07465_(_00698_, _00697_, _00641_);
    and _07466_(_00699_, _00698_, _00695_);
    or _07467_(_00700_, _00620_, _00582_);
    xor _07468_(_00701_, _00582_, _00128_);
    or _07469_(_00702_, _00701_, _00641_);
    and _07470_(_00703_, _00702_, _00700_);
    nand _07471_(_00704_, _00703_, _00699_);
    nor _07472_(_00705_, _00704_, _00694_);
    and _07473_(_00706_, _00705_, _05942_);
    and _07474_(_00707_, _00706_, _00682_);
    and _07475_(_00708_, _00229_, _00226_);
    and _07476_(_00709_, _00708_, _05956_);
    nand _07477_(_00710_, _00709_, _00707_);
    or _07478_(_00711_, _00630_, modulus[6]);
    or _07479_(_00712_, _00678_, modulus[5]);
    or _07480_(_00713_, _00712_, _00674_);
    and _07481_(_00714_, _00713_, _00711_);
    or _07482_(_00715_, _00665_, modulus[4]);
    or _07483_(_00716_, _00670_, modulus[3]);
    or _07484_(_00717_, _00716_, _00666_);
    and _07485_(_00718_, _00717_, _00715_);
    or _07486_(_00719_, _00718_, _00680_);
    and _07487_(_00720_, _00719_, _00714_);
    or _07488_(_00721_, _00638_, modulus[2]);
    or _07489_(_00722_, _00644_, modulus[1]);
    or _07490_(_00723_, _00722_, _00639_);
    and _07491_(_00724_, _00723_, _00721_);
    or _07492_(_00725_, _00651_, modulus[0]);
    or _07493_(_00726_, _00656_, _00652_);
    and _07494_(_00727_, _00726_, _00725_);
    or _07495_(_00728_, _00727_, _00646_);
    and _07496_(_00729_, _00728_, _00724_);
    or _07497_(_00730_, _00729_, _00681_);
    and _07498_(_00731_, _00730_, _00720_);
    and _07499_(_00732_, _00693_, _00689_);
    and _07500_(_00733_, _00703_, _00699_);
    or _07501_(_00734_, _00733_, _00694_);
    and _07502_(_00735_, _00734_, _00732_);
    nand _07503_(_00736_, _00705_, _00372_);
    and _07504_(_00737_, _00736_, _00735_);
    not _07505_(_00738_, _00737_);
    nand _07506_(_00739_, _00738_, _00682_);
    nand _07507_(_00740_, _00739_, _00731_);
    and _07508_(_00741_, _00740_, _00708_);
    nand _07509_(_00742_, _00741_, _05956_);
    nand _07510_(_00743_, _00742_, _00710_);
    or _07511_(_00744_, _00743_, _00630_);
    or _07512_(_00745_, _00737_, _00659_);
    and _07513_(_00746_, _00745_, _00729_);
    or _07514_(_00747_, _00746_, _00672_);
    and _07515_(_00748_, _00747_, _00718_);
    or _07516_(_00749_, _00748_, _00679_);
    and _07517_(_00750_, _00749_, _00712_);
    xor _07518_(_00751_, _00750_, _00674_);
    nand _07519_(_00752_, _00751_, _00743_);
    and _07520_(_00753_, _00752_, _00744_);
    and _07521_(_00754_, _00347_, _00346_);
    or _07522_(_00755_, _00743_, _00638_);
    and _07523_(_00756_, _00742_, _00710_);
    or _07524_(_00757_, _00737_, _00658_);
    and _07525_(_00758_, _00757_, _00727_);
    or _07526_(_00759_, _00758_, _00645_);
    and _07527_(_00760_, _00759_, _00722_);
    xnor _07528_(_00761_, _00760_, _00639_);
    or _07529_(_00762_, _00761_, _00756_);
    and _07530_(_00763_, _00762_, _00755_);
    xor _07531_(_00764_, _00763_, _00309_);
    or _07532_(_00765_, _00743_, _00644_);
    xnor _07533_(_00766_, _00758_, _00645_);
    or _07534_(_00767_, _00766_, _00756_);
    and _07535_(_00768_, _00767_, _00765_);
    xor _07536_(_00769_, _00768_, _00183_);
    or _07537_(_00770_, _00769_, _00764_);
    or _07538_(_00771_, _00743_, _00651_);
    and _07539_(_00772_, _00737_, _00656_);
    xnor _07540_(_00773_, _00772_, _00652_);
    or _07541_(_00774_, _00773_, _00756_);
    and _07542_(_00775_, _00774_, _00771_);
    xor _07543_(_00776_, _00775_, _06035_);
    or _07544_(_00777_, _00743_, _00656_);
    xor _07545_(_00778_, _00737_, _00656_);
    or _07546_(_00779_, _00778_, _00756_);
    and _07547_(_00780_, _00779_, _00777_);
    xor _07548_(_00781_, _00780_, _05927_);
    or _07549_(_00782_, _00781_, _00776_);
    or _07550_(_00783_, _00782_, _00770_);
    or _07551_(_00784_, _00743_, _00665_);
    or _07552_(_00785_, _00746_, _00671_);
    and _07553_(_00786_, _00785_, _00716_);
    xnor _07554_(_00787_, _00786_, _00666_);
    or _07555_(_00788_, _00787_, _00756_);
    and _07556_(_00789_, _00788_, _00784_);
    xor _07557_(_00790_, _00789_, _00550_);
    or _07558_(_00791_, _00743_, _00670_);
    xnor _07559_(_00792_, _00746_, _00671_);
    or _07560_(_00793_, _00792_, _00756_);
    and _07561_(_00794_, _00793_, _00791_);
    xor _07562_(_00795_, _00794_, _00429_);
    or _07563_(_00796_, _00795_, _00790_);
    not _07564_(_00797_, modulus[7]);
    xor _07565_(_00798_, _00753_, _00797_);
    or _07566_(_00799_, _00743_, _00678_);
    xnor _07567_(_00800_, _00748_, _00679_);
    or _07568_(_00801_, _00800_, _00756_);
    and _07569_(_00802_, _00801_, _00799_);
    xor _07570_(_00803_, _00802_, _00673_);
    or _07571_(_00804_, _00803_, _00798_);
    or _07572_(_00805_, _00804_, _00796_);
    nor _07573_(_00806_, _00805_, _00783_);
    or _07574_(_00807_, _00743_, _00689_);
    or _07575_(_00808_, _00704_, _00128_);
    and _07576_(_00809_, _00808_, _00733_);
    and _07577_(_00810_, _00809_, _00693_);
    xor _07578_(_00811_, _00810_, _00689_);
    or _07579_(_00812_, _00811_, _00756_);
    and _07580_(_00813_, _00812_, _00807_);
    or _07581_(_00814_, _00743_, _00693_);
    xor _07582_(_00815_, _00809_, _00693_);
    or _07583_(_00816_, _00815_, _00756_);
    and _07584_(_00817_, _00816_, _00814_);
    nand _07585_(_00818_, _00817_, _00813_);
    or _07586_(_00819_, _00743_, _00699_);
    and _07587_(_00820_, _00703_, _00128_);
    xor _07588_(_00821_, _00820_, _00699_);
    or _07589_(_00822_, _00821_, _00756_);
    and _07590_(_00823_, _00822_, _00819_);
    or _07591_(_00824_, _00743_, _00703_);
    xor _07592_(_00825_, _00703_, _00128_);
    or _07593_(_00826_, _00825_, _00756_);
    and _07594_(_00827_, _00826_, _00824_);
    nand _07595_(_00828_, _00827_, _00823_);
    nor _07596_(_00829_, _00828_, _00818_);
    and _07597_(_00830_, _00829_, _05942_);
    and _07598_(_00831_, _00830_, _00806_);
    nand _07599_(_00832_, _00831_, _00754_);
    or _07600_(_00833_, _00753_, modulus[7]);
    or _07601_(_00834_, _00802_, modulus[6]);
    or _07602_(_00835_, _00834_, _00798_);
    and _07603_(_00836_, _00835_, _00833_);
    or _07604_(_00837_, _00789_, modulus[5]);
    or _07605_(_00838_, _00794_, modulus[4]);
    or _07606_(_00839_, _00838_, _00790_);
    and _07607_(_00840_, _00839_, _00837_);
    or _07608_(_00841_, _00840_, _00804_);
    and _07609_(_00842_, _00841_, _00836_);
    or _07610_(_00843_, _00763_, modulus[3]);
    or _07611_(_00844_, _00768_, modulus[2]);
    or _07612_(_00845_, _00844_, _00764_);
    and _07613_(_00846_, _00845_, _00843_);
    or _07614_(_00847_, _00775_, modulus[1]);
    or _07615_(_00848_, _00780_, modulus[0]);
    or _07616_(_00849_, _00848_, _00776_);
    and _07617_(_00850_, _00849_, _00847_);
    or _07618_(_00851_, _00850_, _00770_);
    and _07619_(_00852_, _00851_, _00846_);
    or _07620_(_00853_, _00852_, _00805_);
    and _07621_(_00854_, _00853_, _00842_);
    and _07622_(_00855_, _00817_, _00813_);
    and _07623_(_00856_, _00827_, _00823_);
    or _07624_(_00857_, _00856_, _00818_);
    and _07625_(_00858_, _00857_, _00855_);
    nand _07626_(_00859_, _00829_, _00372_);
    and _07627_(_00860_, _00859_, _00858_);
    not _07628_(_00861_, _00860_);
    nand _07629_(_00862_, _00861_, _00806_);
    nand _07630_(_00863_, _00862_, _00854_);
    nand _07631_(_00864_, _00863_, _00754_);
    nand _07632_(_00865_, _00864_, _00832_);
    or _07633_(_00866_, _00865_, _00753_);
    or _07634_(_00867_, _00860_, _00783_);
    and _07635_(_00868_, _00867_, _00852_);
    or _07636_(_00869_, _00868_, _00796_);
    and _07637_(_00870_, _00869_, _00840_);
    or _07638_(_00871_, _00870_, _00803_);
    and _07639_(_00872_, _00871_, _00834_);
    xor _07640_(_00873_, _00872_, _00798_);
    nand _07641_(_00874_, _00873_, _00865_);
    and _07642_(_00875_, _00874_, _00866_);
    or _07643_(_00876_, _00865_, _00763_);
    or _07644_(_00877_, _00860_, _00782_);
    and _07645_(_00878_, _00877_, _00850_);
    or _07646_(_00879_, _00878_, _00769_);
    and _07647_(_00880_, _00879_, _00844_);
    xor _07648_(_00881_, _00880_, _00764_);
    nand _07649_(_00882_, _00881_, _00865_);
    and _07650_(_00883_, _00882_, _00876_);
    xor _07651_(_00884_, _00883_, _00429_);
    or _07652_(_00885_, _00865_, _00768_);
    and _07653_(_00886_, _00864_, _00832_);
    xnor _07654_(_00887_, _00878_, _00769_);
    or _07655_(_00888_, _00887_, _00886_);
    and _07656_(_00889_, _00888_, _00885_);
    xor _07657_(_00890_, _00889_, _00309_);
    or _07658_(_00891_, _00890_, _00884_);
    or _07659_(_00892_, _00865_, _00775_);
    or _07660_(_00893_, _00860_, _00781_);
    and _07661_(_00894_, _00893_, _00848_);
    xnor _07662_(_00895_, _00894_, _00776_);
    or _07663_(_00896_, _00895_, _00886_);
    and _07664_(_00897_, _00896_, _00892_);
    xor _07665_(_00898_, _00897_, _00183_);
    or _07666_(_00899_, _00865_, _00780_);
    xnor _07667_(_00900_, _00860_, _00781_);
    or _07668_(_00901_, _00900_, _00886_);
    and _07669_(_00902_, _00901_, _00899_);
    xor _07670_(_00903_, _00902_, _06035_);
    or _07671_(_00904_, _00903_, _00898_);
    or _07672_(_00905_, _00904_, _00891_);
    or _07673_(_00906_, _00865_, _00789_);
    or _07674_(_00907_, _00868_, _00795_);
    and _07675_(_00908_, _00907_, _00838_);
    xor _07676_(_00909_, _00908_, _00790_);
    nand _07677_(_00910_, _00909_, _00865_);
    and _07678_(_00911_, _00910_, _00906_);
    xor _07679_(_00912_, _00911_, _00673_);
    or _07680_(_00913_, _00865_, _00794_);
    xnor _07681_(_00914_, _00868_, _00795_);
    or _07682_(_00915_, _00914_, _00886_);
    and _07683_(_00916_, _00915_, _00913_);
    xor _07684_(_00917_, _00916_, _00550_);
    or _07685_(_00918_, _00917_, _00912_);
    not _07686_(_00919_, modulus[8]);
    xor _07687_(_00920_, _00875_, _00919_);
    or _07688_(_00921_, _00865_, _00802_);
    xor _07689_(_00922_, _00870_, _00803_);
    nand _07690_(_00923_, _00922_, _00865_);
    and _07691_(_00924_, _00923_, _00921_);
    xor _07692_(_00925_, _00924_, _00797_);
    or _07693_(_00926_, _00925_, _00920_);
    or _07694_(_00927_, _00926_, _00918_);
    nor _07695_(_00928_, _00927_, _00905_);
    or _07696_(_00929_, _00865_, _00813_);
    or _07697_(_00930_, _00828_, _00128_);
    and _07698_(_00931_, _00930_, _00856_);
    and _07699_(_00932_, _00931_, _00817_);
    xor _07700_(_00933_, _00932_, _00813_);
    or _07701_(_00934_, _00933_, _00886_);
    and _07702_(_00935_, _00934_, _00929_);
    xor _07703_(_00936_, _00935_, _05927_);
    or _07704_(_00937_, _00865_, _00817_);
    xor _07705_(_00938_, _00931_, _00817_);
    or _07706_(_00939_, _00938_, _00886_);
    and _07707_(_00940_, _00939_, _00937_);
    not _07708_(_00941_, _00940_);
    or _07709_(_00942_, _00941_, _00936_);
    or _07710_(_00943_, _00865_, _00823_);
    and _07711_(_00944_, _00827_, _00128_);
    xor _07712_(_00945_, _00944_, _00823_);
    or _07713_(_00946_, _00945_, _00886_);
    and _07714_(_00947_, _00946_, _00943_);
    or _07715_(_00948_, _00865_, _00827_);
    xor _07716_(_00949_, _00827_, _00128_);
    or _07717_(_00950_, _00949_, _00886_);
    and _07718_(_00951_, _00950_, _00948_);
    nand _07719_(_00952_, _00951_, _00947_);
    nor _07720_(_00953_, _00952_, _00942_);
    and _07721_(_00954_, _00953_, _05942_);
    and _07722_(_00955_, _00954_, _00928_);
    and _07723_(_00956_, _00955_, _05959_);
    not _07724_(_00957_, _00956_);
    or _07725_(_00958_, _00875_, modulus[8]);
    or _07726_(_00959_, _00924_, modulus[7]);
    or _07727_(_00960_, _00959_, _00920_);
    and _07728_(_00961_, _00960_, _00958_);
    or _07729_(_00962_, _00911_, modulus[6]);
    or _07730_(_00963_, _00916_, modulus[5]);
    or _07731_(_00964_, _00963_, _00912_);
    and _07732_(_00965_, _00964_, _00962_);
    or _07733_(_00966_, _00965_, _00926_);
    and _07734_(_00967_, _00966_, _00961_);
    or _07735_(_00968_, _00883_, modulus[4]);
    or _07736_(_00969_, _00889_, modulus[3]);
    or _07737_(_00970_, _00969_, _00884_);
    and _07738_(_00971_, _00970_, _00968_);
    or _07739_(_00972_, _00897_, modulus[2]);
    or _07740_(_00973_, _00902_, modulus[1]);
    or _07741_(_00974_, _00973_, _00898_);
    and _07742_(_00975_, _00974_, _00972_);
    or _07743_(_00976_, _00975_, _00891_);
    and _07744_(_00977_, _00976_, _00971_);
    or _07745_(_00978_, _00977_, _00927_);
    and _07746_(_00979_, _00978_, _00967_);
    or _07747_(_00980_, _00935_, modulus[0]);
    or _07748_(_00981_, _00940_, _00936_);
    and _07749_(_00982_, _00981_, _00980_);
    and _07750_(_00983_, _00951_, _00947_);
    or _07751_(_00984_, _00983_, _00942_);
    and _07752_(_00985_, _00984_, _00982_);
    nand _07753_(_00986_, _00953_, _00372_);
    and _07754_(_00987_, _00986_, _00985_);
    not _07755_(_00988_, _00987_);
    nand _07756_(_00989_, _00988_, _00928_);
    nand _07757_(_00990_, _00989_, _00979_);
    and _07758_(_00991_, _00990_, _05955_);
    and _07759_(_00992_, _00991_, _05957_);
    nand _07760_(_00993_, _00992_, _05956_);
    nand _07761_(_00994_, _00993_, _00957_);
    or _07762_(_00995_, _00994_, _00875_);
    or _07763_(_00996_, _00987_, _00905_);
    and _07764_(_00997_, _00996_, _00977_);
    or _07765_(_00998_, _00997_, _00918_);
    and _07766_(_00999_, _00998_, _00965_);
    or _07767_(_01000_, _00999_, _00925_);
    and _07768_(_01001_, _01000_, _00959_);
    xor _07769_(_01002_, _01001_, _00920_);
    nand _07770_(_01003_, _01002_, _00994_);
    and _07771_(_01004_, _01003_, _00995_);
    or _07772_(_01005_, _00994_, _00883_);
    and _07773_(_01006_, _00993_, _00957_);
    or _07774_(_01007_, _00987_, _00904_);
    and _07775_(_01008_, _01007_, _00975_);
    or _07776_(_01009_, _01008_, _00890_);
    and _07777_(_01010_, _01009_, _00969_);
    xnor _07778_(_01011_, _01010_, _00884_);
    or _07779_(_01012_, _01011_, _01006_);
    and _07780_(_01013_, _01012_, _01005_);
    xor _07781_(_01014_, _01013_, _00550_);
    or _07782_(_01015_, _00994_, _00889_);
    xnor _07783_(_01016_, _01008_, _00890_);
    or _07784_(_01017_, _01016_, _01006_);
    and _07785_(_01018_, _01017_, _01015_);
    xor _07786_(_01019_, _01018_, _00429_);
    or _07787_(_01020_, _01019_, _01014_);
    or _07788_(_01021_, _00994_, _00897_);
    or _07789_(_01022_, _00987_, _00903_);
    and _07790_(_01023_, _01022_, _00973_);
    xnor _07791_(_01024_, _01023_, _00898_);
    or _07792_(_01025_, _01024_, _01006_);
    and _07793_(_01026_, _01025_, _01021_);
    xor _07794_(_01027_, _01026_, _00309_);
    or _07795_(_01028_, _00994_, _00902_);
    xnor _07796_(_01029_, _00987_, _00903_);
    or _07797_(_01030_, _01029_, _01006_);
    and _07798_(_01031_, _01030_, _01028_);
    xor _07799_(_01032_, _01031_, _00183_);
    or _07800_(_01033_, _01032_, _01027_);
    or _07801_(_01034_, _01033_, _01020_);
    or _07802_(_01035_, _00994_, _00911_);
    or _07803_(_01036_, _00997_, _00917_);
    and _07804_(_01037_, _01036_, _00963_);
    xnor _07805_(_01038_, _01037_, _00912_);
    or _07806_(_01039_, _01038_, _01006_);
    and _07807_(_01040_, _01039_, _01035_);
    xor _07808_(_01041_, _01040_, _00797_);
    or _07809_(_01042_, _00994_, _00916_);
    xnor _07810_(_01043_, _00997_, _00917_);
    or _07811_(_01044_, _01043_, _01006_);
    and _07812_(_01045_, _01044_, _01042_);
    xor _07813_(_01046_, _01045_, _00673_);
    or _07814_(_01047_, _01046_, _01041_);
    not _07815_(_01048_, modulus[9]);
    xor _07816_(_01049_, _01004_, _01048_);
    or _07817_(_01050_, _00994_, _00924_);
    xnor _07818_(_01051_, _00999_, _00925_);
    or _07819_(_01052_, _01051_, _01006_);
    and _07820_(_01053_, _01052_, _01050_);
    xor _07821_(_01054_, _01053_, _00919_);
    or _07822_(_01055_, _01054_, _01049_);
    or _07823_(_01056_, _01055_, _01047_);
    nor _07824_(_01057_, _01056_, _01034_);
    or _07825_(_01058_, _00994_, _00935_);
    or _07826_(_01059_, _00952_, _00128_);
    and _07827_(_01060_, _01059_, _00983_);
    and _07828_(_01061_, _01060_, _00940_);
    xnor _07829_(_01062_, _01061_, _00936_);
    or _07830_(_01063_, _01062_, _01006_);
    and _07831_(_01064_, _01063_, _01058_);
    xor _07832_(_01065_, _01064_, _06035_);
    or _07833_(_01066_, _00994_, _00940_);
    xor _07834_(_01067_, _01060_, _00940_);
    or _07835_(_01068_, _01067_, _01006_);
    and _07836_(_01069_, _01068_, _01066_);
    xor _07837_(_01070_, _01069_, _05927_);
    or _07838_(_01071_, _01070_, _01065_);
    or _07839_(_01072_, _00994_, _00947_);
    and _07840_(_01073_, _00951_, _00128_);
    xor _07841_(_01074_, _01073_, _00947_);
    or _07842_(_01075_, _01074_, _01006_);
    and _07843_(_01076_, _01075_, _01072_);
    or _07844_(_01077_, _00994_, _00951_);
    xor _07845_(_01078_, _00951_, _00128_);
    or _07846_(_01079_, _01078_, _01006_);
    and _07847_(_01080_, _01079_, _01077_);
    nand _07848_(_01081_, _01080_, _01076_);
    nor _07849_(_01082_, _01081_, _01071_);
    and _07850_(_01083_, _01082_, _05942_);
    and _07851_(_01084_, _01083_, _01057_);
    and _07852_(_01085_, _01084_, _06075_);
    not _07853_(_01086_, _01085_);
    or _07854_(_01087_, _01004_, modulus[9]);
    or _07855_(_01088_, _01053_, modulus[8]);
    or _07856_(_01089_, _01088_, _01049_);
    and _07857_(_01090_, _01089_, _01087_);
    or _07858_(_01091_, _01040_, modulus[7]);
    or _07859_(_01092_, _01045_, modulus[6]);
    or _07860_(_01093_, _01092_, _01041_);
    and _07861_(_01094_, _01093_, _01091_);
    or _07862_(_01095_, _01094_, _01055_);
    and _07863_(_01096_, _01095_, _01090_);
    or _07864_(_01097_, _01013_, modulus[5]);
    or _07865_(_01098_, _01018_, modulus[4]);
    or _07866_(_01099_, _01098_, _01014_);
    and _07867_(_01100_, _01099_, _01097_);
    or _07868_(_01101_, _01026_, modulus[3]);
    or _07869_(_01102_, _01031_, modulus[2]);
    or _07870_(_01103_, _01102_, _01027_);
    and _07871_(_01104_, _01103_, _01101_);
    or _07872_(_01105_, _01104_, _01020_);
    and _07873_(_01106_, _01105_, _01100_);
    or _07874_(_01107_, _01106_, _01056_);
    and _07875_(_01108_, _01107_, _01096_);
    or _07876_(_01109_, _01064_, modulus[1]);
    or _07877_(_01110_, _01069_, modulus[0]);
    or _07878_(_01111_, _01110_, _01065_);
    and _07879_(_01112_, _01111_, _01109_);
    and _07880_(_01113_, _01080_, _01076_);
    or _07881_(_01114_, _01113_, _01071_);
    and _07882_(_01115_, _01114_, _01112_);
    nand _07883_(_01116_, _01082_, _00372_);
    and _07884_(_01117_, _01116_, _01115_);
    not _07885_(_01118_, _01117_);
    nand _07886_(_01119_, _01118_, _01057_);
    nand _07887_(_01120_, _01119_, _01108_);
    and _07888_(_01121_, _01120_, _06074_);
    nand _07889_(_01122_, _01121_, _06071_);
    nand _07890_(_01123_, _01122_, _01086_);
    or _07891_(_01124_, _01123_, _01004_);
    or _07892_(_01125_, _01117_, _01034_);
    and _07893_(_01126_, _01125_, _01106_);
    or _07894_(_01127_, _01126_, _01047_);
    and _07895_(_01128_, _01127_, _01094_);
    or _07896_(_01129_, _01128_, _01054_);
    and _07897_(_01130_, _01129_, _01088_);
    xor _07898_(_01131_, _01130_, _01049_);
    nand _07899_(_01132_, _01131_, _01123_);
    and _07900_(_01133_, _01132_, _01124_);
    or _07901_(_01134_, _01123_, _01013_);
    or _07902_(_01135_, _01117_, _01033_);
    and _07903_(_01136_, _01135_, _01104_);
    or _07904_(_01137_, _01136_, _01019_);
    and _07905_(_01139_, _01137_, _01098_);
    xor _07906_(_01140_, _01139_, _01014_);
    nand _07907_(_01141_, _01140_, _01123_);
    and _07908_(_01142_, _01141_, _01134_);
    xor _07909_(_01143_, _01142_, _00673_);
    or _07910_(_01144_, _01123_, _01018_);
    and _07911_(_01145_, _01122_, _01086_);
    xnor _07912_(_01146_, _01136_, _01019_);
    or _07913_(_01147_, _01146_, _01145_);
    and _07914_(_01148_, _01147_, _01144_);
    xor _07915_(_01150_, _01148_, _00550_);
    or _07916_(_01151_, _01150_, _01143_);
    or _07917_(_01152_, _01123_, _01026_);
    or _07918_(_01153_, _01117_, _01032_);
    and _07919_(_01154_, _01153_, _01102_);
    xnor _07920_(_01155_, _01154_, _01027_);
    or _07921_(_01156_, _01155_, _01145_);
    and _07922_(_01157_, _01156_, _01152_);
    xor _07923_(_01158_, _01157_, _00429_);
    or _07924_(_01159_, _01123_, _01031_);
    xnor _07925_(_01161_, _01117_, _01032_);
    or _07926_(_01162_, _01161_, _01145_);
    and _07927_(_01163_, _01162_, _01159_);
    xor _07928_(_01164_, _01163_, _00309_);
    or _07929_(_01165_, _01164_, _01158_);
    or _07930_(_01166_, _01165_, _01151_);
    or _07931_(_01167_, _01123_, _01040_);
    or _07932_(_01168_, _01126_, _01046_);
    and _07933_(_01169_, _01168_, _01092_);
    xor _07934_(_01170_, _01169_, _01041_);
    nand _07935_(_01172_, _01170_, _01123_);
    and _07936_(_01173_, _01172_, _01167_);
    xor _07937_(_01174_, _01173_, _00919_);
    or _07938_(_01175_, _01123_, _01045_);
    xnor _07939_(_01176_, _01126_, _01046_);
    or _07940_(_01177_, _01176_, _01145_);
    and _07941_(_01178_, _01177_, _01175_);
    xor _07942_(_01179_, _01178_, _00797_);
    or _07943_(_01180_, _01179_, _01174_);
    not _07944_(_01181_, modulus[10]);
    xor _07945_(_01183_, _01133_, _01181_);
    or _07946_(_01184_, _01123_, _01053_);
    xor _07947_(_01185_, _01128_, _01054_);
    nand _07948_(_01186_, _01185_, _01123_);
    and _07949_(_01187_, _01186_, _01184_);
    xor _07950_(_01188_, _01187_, _01048_);
    or _07951_(_01189_, _01188_, _01183_);
    or _07952_(_01190_, _01189_, _01180_);
    nor _07953_(_01191_, _01190_, _01166_);
    or _07954_(_01192_, _01123_, _01064_);
    or _07955_(_01194_, _01081_, _00128_);
    and _07956_(_01195_, _01194_, _01113_);
    or _07957_(_01196_, _01195_, _01070_);
    and _07958_(_01197_, _01196_, _01110_);
    xnor _07959_(_01198_, _01197_, _01065_);
    or _07960_(_01199_, _01198_, _01145_);
    and _07961_(_01200_, _01199_, _01192_);
    xor _07962_(_01201_, _01200_, _00183_);
    or _07963_(_01202_, _01123_, _01069_);
    xnor _07964_(_01203_, _01195_, _01070_);
    or _07965_(_01205_, _01203_, _01145_);
    and _07966_(_01206_, _01205_, _01202_);
    xor _07967_(_01207_, _01206_, _06035_);
    or _07968_(_01208_, _01207_, _01201_);
    or _07969_(_01209_, _01123_, _01076_);
    and _07970_(_01210_, _01080_, _00128_);
    xor _07971_(_01211_, _01210_, _01076_);
    or _07972_(_01212_, _01211_, _01145_);
    and _07973_(_01213_, _01212_, _01209_);
    xor _07974_(_01214_, _01213_, _05927_);
    or _07975_(_01216_, _01123_, _01080_);
    xor _07976_(_01217_, _01080_, _00128_);
    or _07977_(_01218_, _01217_, _01145_);
    and _07978_(_01219_, _01218_, _01216_);
    not _07979_(_01220_, _01219_);
    or _07980_(_01221_, _01220_, _01214_);
    nor _07981_(_01222_, _01221_, _01208_);
    and _07982_(_01223_, _01222_, _05942_);
    and _07983_(_01224_, _01223_, _01191_);
    nand _07984_(_01225_, _01224_, _00230_);
    or _07985_(_01227_, _01133_, modulus[10]);
    or _07986_(_01228_, _01187_, modulus[9]);
    or _07987_(_01229_, _01228_, _01183_);
    and _07988_(_01230_, _01229_, _01227_);
    or _07989_(_01231_, _01173_, modulus[8]);
    or _07990_(_01232_, _01178_, modulus[7]);
    or _07991_(_01233_, _01232_, _01174_);
    and _07992_(_01234_, _01233_, _01231_);
    or _07993_(_01235_, _01234_, _01189_);
    and _07994_(_01236_, _01235_, _01230_);
    or _07995_(_01238_, _01142_, modulus[6]);
    or _07996_(_01239_, _01148_, modulus[5]);
    or _07997_(_01240_, _01239_, _01143_);
    and _07998_(_01241_, _01240_, _01238_);
    or _07999_(_01242_, _01157_, modulus[4]);
    or _08000_(_01243_, _01163_, modulus[3]);
    or _08001_(_01244_, _01243_, _01158_);
    and _08002_(_01245_, _01244_, _01242_);
    or _08003_(_01246_, _01245_, _01151_);
    and _08004_(_01247_, _01246_, _01241_);
    or _08005_(_01249_, _01247_, _01190_);
    and _08006_(_01250_, _01249_, _01236_);
    or _08007_(_01251_, _01200_, modulus[2]);
    or _08008_(_01252_, _01206_, modulus[1]);
    or _08009_(_01253_, _01252_, _01201_);
    and _08010_(_01254_, _01253_, _01251_);
    or _08011_(_01255_, _01213_, modulus[0]);
    or _08012_(_01256_, _01219_, _01214_);
    and _08013_(_01257_, _01256_, _01255_);
    or _08014_(_01258_, _01257_, _01208_);
    and _08015_(_01260_, _01258_, _01254_);
    nand _08016_(_01261_, _01222_, _00372_);
    nand _08017_(_01262_, _01261_, _01260_);
    nand _08018_(_01263_, _01262_, _01191_);
    nand _08019_(_01264_, _01263_, _01250_);
    and _08020_(_01265_, _01264_, _00229_);
    nand _08021_(_01266_, _01265_, _05956_);
    nand _08022_(_01267_, _01266_, _01225_);
    or _08023_(_01268_, _01267_, _01133_);
    not _08024_(_01269_, _01262_);
    or _08025_(_01271_, _01269_, _01166_);
    and _08026_(_01272_, _01271_, _01247_);
    or _08027_(_01273_, _01272_, _01180_);
    and _08028_(_01274_, _01273_, _01234_);
    or _08029_(_01275_, _01274_, _01188_);
    and _08030_(_01276_, _01275_, _01228_);
    xor _08031_(_01277_, _01276_, _01183_);
    nand _08032_(_01278_, _01277_, _01267_);
    and _08033_(_01279_, _01278_, _01268_);
    or _08034_(_01280_, _01267_, _01142_);
    or _08035_(_01282_, _01269_, _01165_);
    and _08036_(_01283_, _01282_, _01245_);
    or _08037_(_01284_, _01283_, _01150_);
    and _08038_(_01285_, _01284_, _01239_);
    xor _08039_(_01286_, _01285_, _01143_);
    nand _08040_(_01287_, _01286_, _01267_);
    and _08041_(_01288_, _01287_, _01280_);
    xor _08042_(_01289_, _01288_, _00797_);
    or _08043_(_01290_, _01267_, _01148_);
    and _08044_(_01291_, _01266_, _01225_);
    xnor _08045_(_01293_, _01283_, _01150_);
    or _08046_(_01294_, _01293_, _01291_);
    and _08047_(_01295_, _01294_, _01290_);
    xor _08048_(_01296_, _01295_, _00673_);
    or _08049_(_01297_, _01296_, _01289_);
    or _08050_(_01298_, _01267_, _01157_);
    or _08051_(_01299_, _01269_, _01164_);
    and _08052_(_01300_, _01299_, _01243_);
    xnor _08053_(_01301_, _01300_, _01158_);
    or _08054_(_01302_, _01301_, _01291_);
    and _08055_(_01304_, _01302_, _01298_);
    xor _08056_(_01305_, _01304_, _00550_);
    or _08057_(_01306_, _01267_, _01163_);
    xor _08058_(_01307_, _01262_, _01164_);
    or _08059_(_01308_, _01307_, _01291_);
    and _08060_(_01309_, _01308_, _01306_);
    xor _08061_(_01310_, _01309_, _00429_);
    or _08062_(_01311_, _01310_, _01305_);
    or _08063_(_01312_, _01311_, _01297_);
    or _08064_(_01313_, _01267_, _01173_);
    or _08065_(_01315_, _01272_, _01179_);
    and _08066_(_01316_, _01315_, _01232_);
    xor _08067_(_01317_, _01316_, _01174_);
    nand _08068_(_01318_, _01317_, _01267_);
    and _08069_(_01319_, _01318_, _01313_);
    xor _08070_(_01320_, _01319_, _01048_);
    or _08071_(_01321_, _01267_, _01178_);
    xnor _08072_(_01322_, _01272_, _01179_);
    or _08073_(_01323_, _01322_, _01291_);
    and _08074_(_01324_, _01323_, _01321_);
    xor _08075_(_01326_, _01324_, _00919_);
    or _08076_(_01327_, _01326_, _01320_);
    not _08077_(_01328_, modulus[11]);
    xor _08078_(_01329_, _01279_, _01328_);
    or _08079_(_01330_, _01267_, _01187_);
    xor _08080_(_01331_, _01274_, _01188_);
    nand _08081_(_01332_, _01331_, _01267_);
    and _08082_(_01333_, _01332_, _01330_);
    xor _08083_(_01334_, _01333_, _01181_);
    or _08084_(_01335_, _01334_, _01329_);
    or _08085_(_01337_, _01335_, _01327_);
    nor _08086_(_01338_, _01337_, _01312_);
    or _08087_(_01339_, _01267_, _01200_);
    or _08088_(_01340_, _01221_, _00128_);
    and _08089_(_01341_, _01340_, _01257_);
    or _08090_(_01342_, _01341_, _01207_);
    and _08091_(_01343_, _01342_, _01252_);
    xnor _08092_(_01344_, _01343_, _01201_);
    or _08093_(_01345_, _01344_, _01291_);
    and _08094_(_01346_, _01345_, _01339_);
    xor _08095_(_01348_, _01346_, _00309_);
    or _08096_(_01349_, _01267_, _01206_);
    xnor _08097_(_01350_, _01341_, _01207_);
    or _08098_(_01351_, _01350_, _01291_);
    and _08099_(_01352_, _01351_, _01349_);
    xor _08100_(_01353_, _01352_, _00183_);
    or _08101_(_01354_, _01353_, _01348_);
    or _08102_(_01355_, _01267_, _01213_);
    and _08103_(_01356_, _01219_, _00128_);
    xnor _08104_(_01357_, _01356_, _01214_);
    or _08105_(_01359_, _01357_, _01291_);
    and _08106_(_01360_, _01359_, _01355_);
    xor _08107_(_01361_, _01360_, _06035_);
    or _08108_(_01362_, _01267_, _01219_);
    xor _08109_(_01363_, _01219_, _00128_);
    or _08110_(_01364_, _01363_, _01291_);
    and _08111_(_01365_, _01364_, _01362_);
    xor _08112_(_01366_, _01365_, _05927_);
    or _08113_(_01367_, _01366_, _01361_);
    nor _08114_(_01368_, _01367_, _01354_);
    and _08115_(_01370_, _01368_, _05942_);
    and _08116_(_01371_, _01370_, _01338_);
    nand _08117_(_01372_, _01371_, _00346_);
    or _08118_(_01373_, _01279_, modulus[11]);
    or _08119_(_01374_, _01333_, modulus[10]);
    or _08120_(_01375_, _01374_, _01329_);
    and _08121_(_01376_, _01375_, _01373_);
    or _08122_(_01377_, _01319_, modulus[9]);
    or _08123_(_01378_, _01324_, modulus[8]);
    or _08124_(_01379_, _01378_, _01320_);
    and _08125_(_01381_, _01379_, _01377_);
    or _08126_(_01382_, _01381_, _01335_);
    and _08127_(_01383_, _01382_, _01376_);
    or _08128_(_01384_, _01288_, modulus[7]);
    or _08129_(_01385_, _01295_, modulus[6]);
    or _08130_(_01386_, _01385_, _01289_);
    and _08131_(_01387_, _01386_, _01384_);
    or _08132_(_01388_, _01304_, modulus[5]);
    or _08133_(_01389_, _01309_, modulus[4]);
    or _08134_(_01390_, _01389_, _01305_);
    and _08135_(_01392_, _01390_, _01388_);
    or _08136_(_01393_, _01392_, _01297_);
    and _08137_(_01394_, _01393_, _01387_);
    or _08138_(_01395_, _01394_, _01337_);
    and _08139_(_01396_, _01395_, _01383_);
    or _08140_(_01397_, _01346_, modulus[3]);
    or _08141_(_01398_, _01352_, modulus[2]);
    or _08142_(_01399_, _01398_, _01348_);
    and _08143_(_01400_, _01399_, _01397_);
    or _08144_(_01401_, _01360_, modulus[1]);
    or _08145_(_01403_, _01365_, modulus[0]);
    or _08146_(_01404_, _01403_, _01361_);
    and _08147_(_01405_, _01404_, _01401_);
    or _08148_(_01406_, _01405_, _01354_);
    and _08149_(_01407_, _01406_, _01400_);
    nand _08150_(_01408_, _01368_, _00372_);
    and _08151_(_01409_, _01408_, _01407_);
    not _08152_(_01410_, _01409_);
    nand _08153_(_01411_, _01410_, _01338_);
    nand _08154_(_01412_, _01411_, _01396_);
    nand _08155_(_01414_, _01412_, _00346_);
    nand _08156_(_01415_, _01414_, _01372_);
    or _08157_(_01416_, _01415_, _01279_);
    or _08158_(_01417_, _01409_, _01312_);
    and _08159_(_01418_, _01417_, _01394_);
    or _08160_(_01419_, _01418_, _01327_);
    and _08161_(_01420_, _01419_, _01381_);
    or _08162_(_01421_, _01420_, _01334_);
    and _08163_(_01422_, _01421_, _01374_);
    xor _08164_(_01423_, _01422_, _01329_);
    nand _08165_(_01425_, _01423_, _01415_);
    and _08166_(_01426_, _01425_, _01416_);
    or _08167_(_01427_, _01415_, _01288_);
    or _08168_(_01428_, _01409_, _01311_);
    and _08169_(_01429_, _01428_, _01392_);
    or _08170_(_01430_, _01429_, _01296_);
    and _08171_(_01431_, _01430_, _01385_);
    xor _08172_(_01432_, _01431_, _01289_);
    nand _08173_(_01433_, _01432_, _01415_);
    and _08174_(_01434_, _01433_, _01427_);
    xor _08175_(_01436_, _01434_, _00919_);
    or _08176_(_01437_, _01415_, _01295_);
    xor _08177_(_01438_, _01429_, _01296_);
    nand _08178_(_01439_, _01438_, _01415_);
    and _08179_(_01440_, _01439_, _01437_);
    xor _08180_(_01441_, _01440_, _00797_);
    or _08181_(_01442_, _01441_, _01436_);
    or _08182_(_01443_, _01415_, _01304_);
    or _08183_(_01444_, _01409_, _01310_);
    and _08184_(_01445_, _01444_, _01389_);
    xor _08185_(_01447_, _01445_, _01305_);
    nand _08186_(_01448_, _01447_, _01415_);
    and _08187_(_01449_, _01448_, _01443_);
    xor _08188_(_01450_, _01449_, _00673_);
    or _08189_(_01451_, _01415_, _01309_);
    and _08190_(_01452_, _01414_, _01372_);
    xnor _08191_(_01453_, _01409_, _01310_);
    or _08192_(_01454_, _01453_, _01452_);
    and _08193_(_01455_, _01454_, _01451_);
    xor _08194_(_01456_, _01455_, _00550_);
    or _08195_(_01458_, _01456_, _01450_);
    or _08196_(_01459_, _01458_, _01442_);
    or _08197_(_01460_, _01415_, _01319_);
    or _08198_(_01461_, _01418_, _01326_);
    and _08199_(_01462_, _01461_, _01378_);
    xor _08200_(_01463_, _01462_, _01320_);
    nand _08201_(_01464_, _01463_, _01415_);
    and _08202_(_01465_, _01464_, _01460_);
    xor _08203_(_01466_, _01465_, _01181_);
    or _08204_(_01467_, _01415_, _01324_);
    xor _08205_(_01469_, _01418_, _01326_);
    nand _08206_(_01470_, _01469_, _01415_);
    and _08207_(_01471_, _01470_, _01467_);
    xor _08208_(_01472_, _01471_, _01048_);
    or _08209_(_01473_, _01472_, _01466_);
    not _08210_(_01474_, modulus[12]);
    xor _08211_(_01475_, _01426_, _01474_);
    or _08212_(_01476_, _01415_, _01333_);
    xor _08213_(_01477_, _01420_, _01334_);
    nand _08214_(_01478_, _01477_, _01415_);
    and _08215_(_01480_, _01478_, _01476_);
    xor _08216_(_01481_, _01480_, _01328_);
    or _08217_(_01482_, _01481_, _01475_);
    or _08218_(_01483_, _01482_, _01473_);
    or _08219_(_01484_, _01483_, _01459_);
    or _08220_(_01485_, _01415_, _01346_);
    or _08221_(_01486_, _01367_, _00128_);
    and _08222_(_01487_, _01486_, _01405_);
    or _08223_(_01488_, _01487_, _01353_);
    and _08224_(_01489_, _01488_, _01398_);
    xnor _08225_(_01491_, _01489_, _01348_);
    or _08226_(_01492_, _01491_, _01452_);
    and _08227_(_01493_, _01492_, _01485_);
    xor _08228_(_01494_, _01493_, _00429_);
    or _08229_(_01495_, _01415_, _01352_);
    xnor _08230_(_01496_, _01487_, _01353_);
    or _08231_(_01497_, _01496_, _01452_);
    and _08232_(_01498_, _01497_, _01495_);
    xor _08233_(_01499_, _01498_, _00309_);
    or _08234_(_01500_, _01499_, _01494_);
    or _08235_(_01502_, _01415_, _01360_);
    or _08236_(_01503_, _01366_, _00128_);
    and _08237_(_01504_, _01503_, _01403_);
    xnor _08238_(_01505_, _01504_, _01361_);
    or _08239_(_01506_, _01505_, _01452_);
    and _08240_(_01507_, _01506_, _01502_);
    xor _08241_(_01508_, _01507_, _00183_);
    or _08242_(_01509_, _01415_, _01365_);
    xor _08243_(_01510_, _01366_, _00372_);
    or _08244_(_01511_, _01510_, _01452_);
    and _08245_(_01513_, _01511_, _01509_);
    xor _08246_(_01514_, _01513_, _06035_);
    or _08247_(_01515_, _01514_, _01508_);
    or _08248_(_01516_, _01515_, _01500_);
    xor _08249_(_01517_, _05980_, modulus[0]);
    and _08250_(_01518_, _01517_, _05981_);
    and _08251_(_01519_, _01518_, _01138_);
    not _08252_(_01520_, _01519_);
    nor _08253_(_01521_, _01520_, _01516_);
    not _08254_(_01522_, _01521_);
    nor _08255_(_01524_, _01522_, _01484_);
    nand _08256_(_01525_, _01524_, _05958_);
    or _08257_(_01526_, _01426_, modulus[12]);
    or _08258_(_01527_, _01480_, modulus[11]);
    or _08259_(_01528_, _01527_, _01475_);
    and _08260_(_01529_, _01528_, _01526_);
    or _08261_(_01530_, _01465_, modulus[10]);
    or _08262_(_01531_, _01471_, modulus[9]);
    or _08263_(_01532_, _01531_, _01466_);
    and _08264_(_01533_, _01532_, _01530_);
    or _08265_(_01535_, _01533_, _01482_);
    and _08266_(_01536_, _01535_, _01529_);
    or _08267_(_01537_, _01434_, modulus[8]);
    or _08268_(_01538_, _01440_, modulus[7]);
    or _08269_(_01539_, _01538_, _01436_);
    and _08270_(_01540_, _01539_, _01537_);
    or _08271_(_01541_, _01449_, modulus[6]);
    or _08272_(_01542_, _01455_, modulus[5]);
    or _08273_(_01543_, _01542_, _01450_);
    and _08274_(_01544_, _01543_, _01541_);
    or _08275_(_01546_, _01544_, _01442_);
    and _08276_(_01547_, _01546_, _01540_);
    or _08277_(_01548_, _01547_, _01483_);
    and _08278_(_01549_, _01548_, _01536_);
    or _08279_(_01550_, _01493_, modulus[4]);
    or _08280_(_01551_, _01498_, modulus[3]);
    or _08281_(_01552_, _01551_, _01494_);
    and _08282_(_01553_, _01552_, _01550_);
    or _08283_(_01554_, _01507_, modulus[2]);
    or _08284_(_01555_, _01513_, modulus[1]);
    or _08285_(_01557_, _01555_, _01508_);
    and _08286_(_01558_, _01557_, _01554_);
    or _08287_(_01559_, _01558_, _01500_);
    and _08288_(_01560_, _01559_, _01553_);
    and _08289_(_01561_, _05980_, modulus[0]);
    or _08290_(_01562_, _01561_, _01516_);
    and _08291_(_01563_, _01562_, _01560_);
    or _08292_(_01564_, _01563_, _01484_);
    nand _08293_(_01565_, _01564_, _01549_);
    and _08294_(_01566_, _01565_, _05957_);
    nand _08295_(_01568_, _01566_, _05956_);
    nand _08296_(_01569_, _01568_, _01525_);
    or _08297_(_01570_, _01569_, _01426_);
    or _08298_(_01571_, _01563_, _01459_);
    and _08299_(_01572_, _01571_, _01547_);
    or _08300_(_01573_, _01572_, _01473_);
    and _08301_(_01574_, _01573_, _01533_);
    or _08302_(_01575_, _01574_, _01481_);
    and _08303_(_01576_, _01575_, _01527_);
    xor _08304_(_01577_, _01576_, _01475_);
    nand _08305_(_01579_, _01577_, _01569_);
    and _08306_(_01580_, _01579_, _01570_);
    or _08307_(_01581_, _01569_, _01434_);
    and _08308_(_01582_, _01568_, _01525_);
    or _08309_(_01583_, _01563_, _01458_);
    and _08310_(_01584_, _01583_, _01544_);
    or _08311_(_01585_, _01584_, _01441_);
    and _08312_(_01586_, _01585_, _01538_);
    xnor _08313_(_01587_, _01586_, _01436_);
    or _08314_(_01588_, _01587_, _01582_);
    and _08315_(_01590_, _01588_, _01581_);
    xor _08316_(_01591_, _01590_, _01048_);
    or _08317_(_01592_, _01569_, _01440_);
    xnor _08318_(_01593_, _01584_, _01441_);
    or _08319_(_01594_, _01593_, _01582_);
    and _08320_(_01595_, _01594_, _01592_);
    xor _08321_(_01596_, _01595_, _00919_);
    or _08322_(_01597_, _01596_, _01591_);
    or _08323_(_01598_, _01569_, _01449_);
    or _08324_(_01599_, _01563_, _01456_);
    and _08325_(_01601_, _01599_, _01542_);
    xnor _08326_(_01602_, _01601_, _01450_);
    or _08327_(_01603_, _01602_, _01582_);
    and _08328_(_01604_, _01603_, _01598_);
    xor _08329_(_01605_, _01604_, _00797_);
    or _08330_(_01606_, _01569_, _01455_);
    xnor _08331_(_01607_, _01563_, _01456_);
    or _08332_(_01608_, _01607_, _01582_);
    and _08333_(_01609_, _01608_, _01606_);
    xor _08334_(_01610_, _01609_, _00673_);
    or _08335_(_01612_, _01610_, _01605_);
    or _08336_(_01613_, _01612_, _01597_);
    or _08337_(_01614_, _01569_, _01465_);
    or _08338_(_01615_, _01572_, _01472_);
    and _08339_(_01616_, _01615_, _01531_);
    xnor _08340_(_01617_, _01616_, _01466_);
    or _08341_(_01618_, _01617_, _01582_);
    and _08342_(_01619_, _01618_, _01614_);
    xor _08343_(_01620_, _01619_, _01328_);
    or _08344_(_01621_, _01569_, _01471_);
    xnor _08345_(_01623_, _01572_, _01472_);
    or _08346_(_01624_, _01623_, _01582_);
    and _08347_(_01625_, _01624_, _01621_);
    xor _08348_(_01626_, _01625_, _01181_);
    or _08349_(_01627_, _01626_, _01620_);
    not _08350_(_01628_, modulus[13]);
    xor _08351_(_01629_, _01580_, _01628_);
    or _08352_(_01630_, _01569_, _01480_);
    xnor _08353_(_01631_, _01574_, _01481_);
    or _08354_(_01632_, _01631_, _01582_);
    and _08355_(_01634_, _01632_, _01630_);
    xor _08356_(_01635_, _01634_, _01474_);
    or _08357_(_01636_, _01635_, _01629_);
    or _08358_(_01637_, _01636_, _01627_);
    nor _08359_(_01638_, _01637_, _01613_);
    or _08360_(_01639_, _01569_, _01493_);
    or _08361_(_01640_, _01561_, _01515_);
    and _08362_(_01641_, _01640_, _01558_);
    or _08363_(_01642_, _01641_, _01499_);
    and _08364_(_01643_, _01642_, _01551_);
    xnor _08365_(_01645_, _01643_, _01494_);
    or _08366_(_01646_, _01645_, _01582_);
    and _08367_(_01647_, _01646_, _01639_);
    xor _08368_(_01648_, _01647_, _00550_);
    or _08369_(_01649_, _01569_, _01498_);
    xnor _08370_(_01650_, _01641_, _01499_);
    or _08371_(_01651_, _01650_, _01582_);
    and _08372_(_01652_, _01651_, _01649_);
    xor _08373_(_01653_, _01652_, _00429_);
    or _08374_(_01654_, _01653_, _01648_);
    or _08375_(_01656_, _01569_, _01507_);
    or _08376_(_01657_, _01561_, _01514_);
    and _08377_(_01658_, _01657_, _01555_);
    xnor _08378_(_01659_, _01658_, _01508_);
    or _08379_(_01660_, _01659_, _01582_);
    and _08380_(_01661_, _01660_, _01656_);
    xor _08381_(_01662_, _01661_, _00309_);
    or _08382_(_01663_, _01569_, _01513_);
    xnor _08383_(_01664_, _01561_, _01514_);
    or _08384_(_01665_, _01664_, _01582_);
    and _08385_(_01667_, _01665_, _01663_);
    xor _08386_(_01668_, _01667_, _00183_);
    or _08387_(_01669_, _01668_, _01662_);
    or _08388_(_01670_, _01669_, _01654_);
    not _08389_(_01671_, _01670_);
    or _08390_(_01672_, _01569_, _05980_);
    or _08391_(_01673_, _01582_, _01517_);
    and _08392_(_01674_, _01673_, _01672_);
    xor _08393_(_01675_, _01674_, _06035_);
    xor _08394_(_01676_, _05981_, _05927_);
    or _08395_(_01677_, _01676_, _01675_);
    nor _08396_(_01678_, _01677_, base[0]);
    and _08397_(_01679_, _01678_, _01671_);
    and _08398_(_01680_, _01679_, _01638_);
    nand _08399_(_01681_, _01680_, _06071_);
    or _08400_(_01682_, _01580_, modulus[13]);
    or _08401_(_01683_, _01634_, modulus[12]);
    or _08402_(_01684_, _01683_, _01629_);
    and _08403_(_01685_, _01684_, _01682_);
    or _08404_(_01686_, _01619_, modulus[11]);
    or _08405_(_01688_, _01625_, modulus[10]);
    or _08406_(_01689_, _01688_, _01620_);
    and _08407_(_01690_, _01689_, _01686_);
    or _08408_(_01691_, _01690_, _01636_);
    and _08409_(_01692_, _01691_, _01685_);
    or _08410_(_01693_, _01590_, modulus[9]);
    or _08411_(_01694_, _01595_, modulus[8]);
    or _08412_(_01695_, _01694_, _01591_);
    and _08413_(_01696_, _01695_, _01693_);
    or _08414_(_01697_, _01604_, modulus[7]);
    or _08415_(_01699_, _01609_, modulus[6]);
    or _08416_(_01700_, _01699_, _01605_);
    and _08417_(_01701_, _01700_, _01697_);
    or _08418_(_01702_, _01701_, _01597_);
    and _08419_(_01703_, _01702_, _01696_);
    or _08420_(_01704_, _01703_, _01637_);
    and _08421_(_01705_, _01704_, _01692_);
    or _08422_(_01706_, _01647_, modulus[5]);
    or _08423_(_01707_, _01652_, modulus[4]);
    or _08424_(_01708_, _01707_, _01648_);
    and _08425_(_01710_, _01708_, _01706_);
    or _08426_(_01711_, _01661_, modulus[3]);
    or _08427_(_01712_, _01667_, modulus[2]);
    or _08428_(_01713_, _01712_, _01662_);
    and _08429_(_01714_, _01713_, _01711_);
    or _08430_(_01715_, _01714_, _01654_);
    and _08431_(_01716_, _01715_, _01710_);
    or _08432_(_01717_, _01674_, modulus[1]);
    or _08433_(_01718_, _05981_, modulus[0]);
    or _08434_(_01719_, _01718_, _01675_);
    and _08435_(_01721_, _01719_, _01717_);
    and _08436_(_01722_, _01721_, _01677_);
    or _08437_(_01723_, _01722_, _01670_);
    and _08438_(_01724_, _01723_, _01716_);
    not _08439_(_01725_, _01724_);
    nand _08440_(_01726_, _01725_, _01638_);
    nand _08441_(_01727_, _01726_, _01705_);
    nand _08442_(_01728_, _01727_, _06071_);
    nand _08443_(_01729_, _01728_, _01681_);
    or _08444_(_01730_, _01729_, _01580_);
    and _08445_(_01732_, _01728_, _01681_);
    or _08446_(_01733_, _01724_, _01613_);
    and _08447_(_01734_, _01733_, _01703_);
    or _08448_(_01735_, _01734_, _01627_);
    and _08449_(_01736_, _01735_, _01690_);
    or _08450_(_01737_, _01736_, _01635_);
    nand _08451_(_01738_, _01737_, _01683_);
    xor _08452_(_01739_, _01738_, _01629_);
    or _08453_(_01740_, _01739_, _01732_);
    and _08454_(_01741_, _01740_, _01730_);
    or _08455_(_01743_, _01729_, _01590_);
    or _08456_(_01744_, _01724_, _01612_);
    and _08457_(_01745_, _01744_, _01701_);
    or _08458_(_01746_, _01745_, _01596_);
    nand _08459_(_01747_, _01746_, _01694_);
    xor _08460_(_01748_, _01747_, _01591_);
    or _08461_(_01749_, _01748_, _01732_);
    and _08462_(_01750_, _01749_, _01743_);
    xor _08463_(_01751_, _01750_, _01181_);
    or _08464_(_01752_, _01729_, _01595_);
    xnor _08465_(_01754_, _01745_, _01596_);
    or _08466_(_01755_, _01754_, _01732_);
    and _08467_(_01756_, _01755_, _01752_);
    xor _08468_(_01757_, _01756_, _01048_);
    or _08469_(_01758_, _01757_, _01751_);
    or _08470_(_01759_, _01729_, _01604_);
    or _08471_(_01760_, _01724_, _01610_);
    nand _08472_(_01761_, _01760_, _01699_);
    xor _08473_(_01762_, _01761_, _01605_);
    or _08474_(_01763_, _01762_, _01732_);
    and _08475_(_01765_, _01763_, _01759_);
    xor _08476_(_01766_, _01765_, _00919_);
    or _08477_(_01767_, _01729_, _01609_);
    xnor _08478_(_01768_, _01724_, _01610_);
    or _08479_(_01769_, _01768_, _01732_);
    and _08480_(_01770_, _01769_, _01767_);
    xor _08481_(_01771_, _01770_, _00797_);
    or _08482_(_01772_, _01771_, _01766_);
    or _08483_(_01773_, _01772_, _01758_);
    or _08484_(_01774_, _01729_, _01619_);
    or _08485_(_01776_, _01734_, _01626_);
    nand _08486_(_01777_, _01776_, _01688_);
    xor _08487_(_01778_, _01777_, _01620_);
    or _08488_(_01779_, _01778_, _01732_);
    and _08489_(_01780_, _01779_, _01774_);
    xor _08490_(_01781_, _01780_, _01474_);
    or _08491_(_01782_, _01729_, _01625_);
    xnor _08492_(_01783_, _01734_, _01626_);
    or _08493_(_01784_, _01783_, _01732_);
    and _08494_(_01785_, _01784_, _01782_);
    xor _08495_(_01787_, _01785_, _01328_);
    or _08496_(_01788_, _01787_, _01781_);
    not _08497_(_01789_, modulus[14]);
    xor _08498_(_01790_, _01741_, _01789_);
    or _08499_(_01791_, _01729_, _01634_);
    xnor _08500_(_01792_, _01736_, _01635_);
    or _08501_(_01793_, _01792_, _01732_);
    and _08502_(_01794_, _01793_, _01791_);
    xor _08503_(_01795_, _01794_, _01628_);
    or _08504_(_01796_, _01795_, _01790_);
    or _08505_(_01798_, _01796_, _01788_);
    or _08506_(_01799_, _01798_, _01773_);
    or _08507_(_01800_, _01729_, _01647_);
    or _08508_(_01801_, _01722_, _01669_);
    and _08509_(_01802_, _01801_, _01714_);
    or _08510_(_01803_, _01802_, _01653_);
    nand _08511_(_01804_, _01803_, _01707_);
    xor _08512_(_01805_, _01804_, _01648_);
    or _08513_(_01806_, _01805_, _01732_);
    and _08514_(_01807_, _01806_, _01800_);
    xor _08515_(_01809_, _01807_, _00673_);
    or _08516_(_01810_, _01729_, _01652_);
    xnor _08517_(_01811_, _01802_, _01653_);
    or _08518_(_01812_, _01811_, _01732_);
    and _08519_(_01813_, _01812_, _01810_);
    xor _08520_(_01814_, _01813_, _00550_);
    or _08521_(_01815_, _01814_, _01809_);
    or _08522_(_01816_, _01729_, _01661_);
    or _08523_(_01817_, _01722_, _01668_);
    nand _08524_(_01818_, _01817_, _01712_);
    xor _08525_(_01820_, _01818_, _01662_);
    or _08526_(_01821_, _01820_, _01732_);
    and _08527_(_01822_, _01821_, _01816_);
    xor _08528_(_01823_, _01822_, _00429_);
    or _08529_(_01824_, _01729_, _01667_);
    xnor _08530_(_01825_, _01722_, _01668_);
    or _08531_(_01826_, _01825_, _01732_);
    and _08532_(_01827_, _01826_, _01824_);
    xor _08533_(_01828_, _01827_, _00309_);
    or _08534_(_01829_, _01828_, _01823_);
    or _08535_(_01831_, _01829_, _01815_);
    or _08536_(_01832_, modulus[0], base[0]);
    or _08537_(_01833_, _01729_, _01674_);
    nand _08538_(_01834_, _05981_, modulus[0]);
    xor _08539_(_01835_, _01834_, _01675_);
    or _08540_(_01836_, _01835_, _01732_);
    and _08541_(_01837_, _01836_, _01833_);
    xor _08542_(_01838_, _01837_, _00183_);
    or _08543_(_01839_, _01729_, _05981_);
    nand _08544_(_01840_, _01729_, _01676_);
    and _08545_(_01842_, _01840_, _01839_);
    xor _08546_(_01843_, _01842_, _06035_);
    or _08547_(_01844_, _01843_, _01838_);
    or _08548_(_01845_, _01844_, _01832_);
    or _08549_(_01846_, _01845_, _01831_);
    nor _08550_(_01847_, _01846_, _01799_);
    or _08551_(_01848_, _01741_, modulus[14]);
    or _08552_(_01849_, _01794_, modulus[13]);
    or _08553_(_01850_, _01849_, _01790_);
    and _08554_(_01851_, _01850_, _01848_);
    or _08555_(_01853_, _01780_, modulus[12]);
    or _08556_(_01854_, _01785_, modulus[11]);
    or _08557_(_01855_, _01854_, _01781_);
    and _08558_(_01856_, _01855_, _01853_);
    or _08559_(_01857_, _01856_, _01796_);
    and _08560_(_01858_, _01857_, _01851_);
    or _08561_(_01859_, _01750_, modulus[10]);
    or _08562_(_01860_, _01756_, modulus[9]);
    or _08563_(_01861_, _01860_, _01751_);
    and _08564_(_01862_, _01861_, _01859_);
    or _08565_(_01864_, _01765_, modulus[8]);
    or _08566_(_01865_, _01770_, modulus[7]);
    or _08567_(_01866_, _01865_, _01766_);
    and _08568_(_01867_, _01866_, _01864_);
    or _08569_(_01868_, _01867_, _01758_);
    and _08570_(_01869_, _01868_, _01862_);
    or _08571_(_01870_, _01869_, _01798_);
    and _08572_(_01871_, _01870_, _01858_);
    or _08573_(_01872_, _01807_, modulus[6]);
    or _08574_(_01873_, _01813_, modulus[5]);
    or _08575_(_01875_, _01873_, _01809_);
    and _08576_(_01876_, _01875_, _01872_);
    or _08577_(_01877_, _01822_, modulus[4]);
    or _08578_(_01878_, _01827_, modulus[3]);
    or _08579_(_01879_, _01878_, _01823_);
    and _08580_(_01880_, _01879_, _01877_);
    or _08581_(_01881_, _01880_, _01815_);
    and _08582_(_01882_, _01881_, _01876_);
    or _08583_(_01883_, _01837_, modulus[2]);
    or _08584_(_01884_, _01842_, modulus[1]);
    or _08585_(_01886_, _01884_, _01838_);
    and _08586_(_01887_, _01886_, _01883_);
    or _08587_(_01888_, _01844_, modulus[0]);
    and _08588_(_01889_, _01888_, _01887_);
    or _08589_(_01890_, _01889_, _01831_);
    and _08590_(_01891_, _01890_, _01882_);
    or _08591_(_01892_, _01891_, _01799_);
    and _08592_(_01893_, _01892_, _01871_);
    or _08593_(_01894_, _01891_, _01773_);
    and _08594_(_01895_, _01894_, _01869_);
    or _08595_(_01897_, _01895_, _01788_);
    and _08596_(_01898_, _01897_, _01856_);
    or _08597_(_01899_, _01898_, _01795_);
    nand _08598_(_01900_, _01899_, _01849_);
    xor _08599_(_01901_, _01900_, _01790_);
    and _08600_(_01902_, _01741_, modulus[15]);
    nand _08601_(_01903_, _01847_, _05956_);
    or _08602_(_01904_, _01893_, modulus[15]);
    nand _08603_(_01905_, _01904_, _01903_);
    or _08604_(_01906_, _01905_, _01741_);
    and _08605_(_01908_, _01904_, _01903_);
    or _08606_(_01909_, _01901_, _01908_);
    and _08607_(_01910_, _01909_, _01906_);
    xor _08608_(_01911_, _01910_, _05956_);
    or _08609_(_01912_, _01905_, _01794_);
    xnor _08610_(_01913_, _01898_, _01795_);
    or _08611_(_01914_, _01913_, _01908_);
    and _08612_(_01915_, _01914_, _01912_);
    nand _08613_(_01916_, _01915_, modulus[14]);
    nor _08614_(_01917_, _01916_, _01911_);
    nor _08615_(_01919_, _01917_, _01902_);
    xor _08616_(_01920_, _01915_, _01789_);
    nor _08617_(_01921_, _01920_, _01911_);
    or _08618_(_01922_, _01905_, _01780_);
    or _08619_(_01923_, _01895_, _01787_);
    nand _08620_(_01924_, _01923_, _01854_);
    xor _08621_(_01925_, _01924_, _01781_);
    or _08622_(_01926_, _01925_, _01908_);
    and _08623_(_01927_, _01926_, _01922_);
    and _08624_(_01928_, _01927_, modulus[13]);
    xor _08625_(_01930_, _01927_, _01628_);
    or _08626_(_01931_, _01905_, _01785_);
    xnor _08627_(_01932_, _01895_, _01787_);
    or _08628_(_01933_, _01932_, _01908_);
    and _08629_(_01934_, _01933_, _01931_);
    nand _08630_(_01935_, _01934_, modulus[12]);
    nor _08631_(_01936_, _01935_, _01930_);
    nor _08632_(_01937_, _01936_, _01928_);
    not _08633_(_01938_, _01937_);
    and _08634_(_01939_, _01938_, _01921_);
    not _08635_(_01941_, _01939_);
    and _08636_(_01942_, _01941_, _01919_);
    xor _08637_(_01943_, _01934_, _01474_);
    nor _08638_(_01944_, _01943_, _01930_);
    and _08639_(_01945_, _01944_, _01921_);
    or _08640_(_01946_, _01905_, _01750_);
    or _08641_(_01947_, _01891_, _01772_);
    and _08642_(_01948_, _01947_, _01867_);
    or _08643_(_01949_, _01948_, _01757_);
    nand _08644_(_01950_, _01949_, _01860_);
    xor _08645_(_01952_, _01950_, _01751_);
    or _08646_(_01953_, _01952_, _01908_);
    and _08647_(_01954_, _01953_, _01946_);
    and _08648_(_01955_, _01954_, modulus[11]);
    xor _08649_(_01956_, _01954_, _01328_);
    or _08650_(_01957_, _01905_, _01756_);
    xnor _08651_(_01958_, _01948_, _01757_);
    or _08652_(_01959_, _01958_, _01908_);
    and _08653_(_01960_, _01959_, _01957_);
    nand _08654_(_01961_, _01960_, modulus[10]);
    nor _08655_(_01963_, _01961_, _01956_);
    nor _08656_(_01964_, _01963_, _01955_);
    xor _08657_(_01965_, _01960_, _01181_);
    or _08658_(_01966_, _01965_, _01956_);
    or _08659_(_01967_, _01905_, _01765_);
    or _08660_(_01968_, _01891_, _01771_);
    nand _08661_(_01969_, _01968_, _01865_);
    xor _08662_(_01970_, _01969_, _01766_);
    or _08663_(_01971_, _01970_, _01908_);
    and _08664_(_01972_, _01971_, _01967_);
    nand _08665_(_01974_, _01972_, modulus[9]);
    xor _08666_(_01975_, _01972_, _01048_);
    or _08667_(_01976_, _01905_, _01770_);
    xnor _08668_(_01977_, _01891_, _01771_);
    or _08669_(_01978_, _01977_, _01908_);
    and _08670_(_01979_, _01978_, _01976_);
    nand _08671_(_01980_, _01979_, modulus[8]);
    or _08672_(_01981_, _01980_, _01975_);
    and _08673_(_01982_, _01981_, _01974_);
    nor _08674_(_01983_, _01982_, _01966_);
    not _08675_(_01985_, _01983_);
    nand _08676_(_01986_, _01985_, _01964_);
    nand _08677_(_01987_, _01986_, _01945_);
    and _08678_(_01988_, _01987_, _01942_);
    xor _08679_(_01989_, _01979_, _00919_);
    or _08680_(_01990_, _01989_, _01975_);
    or _08681_(_01991_, _01990_, _01966_);
    not _08682_(_01992_, _01991_);
    and _08683_(_01993_, _01992_, _01945_);
    or _08684_(_01994_, _01905_, _01807_);
    or _08685_(_01996_, _01889_, _01829_);
    and _08686_(_01997_, _01996_, _01880_);
    or _08687_(_01998_, _01997_, _01814_);
    nand _08688_(_01999_, _01998_, _01873_);
    xor _08689_(_02000_, _01999_, _01809_);
    or _08690_(_02001_, _02000_, _01908_);
    and _08691_(_02002_, _02001_, _01994_);
    and _08692_(_02003_, _02002_, modulus[7]);
    xor _08693_(_02004_, _02002_, _00797_);
    or _08694_(_02005_, _01905_, _01813_);
    xnor _08695_(_02007_, _01997_, _01814_);
    or _08696_(_02008_, _02007_, _01908_);
    and _08697_(_02009_, _02008_, _02005_);
    nand _08698_(_02010_, _02009_, modulus[6]);
    nor _08699_(_02011_, _02010_, _02004_);
    nor _08700_(_02012_, _02011_, _02003_);
    xor _08701_(_02013_, _02009_, _00673_);
    or _08702_(_02014_, _02013_, _02004_);
    or _08703_(_02015_, _01905_, _01822_);
    or _08704_(_02016_, _01889_, _01828_);
    nand _08705_(_02018_, _02016_, _01878_);
    xor _08706_(_02019_, _02018_, _01823_);
    or _08707_(_02020_, _02019_, _01908_);
    and _08708_(_02021_, _02020_, _02015_);
    nand _08709_(_02022_, _02021_, modulus[5]);
    xor _08710_(_02023_, _02021_, _00550_);
    or _08711_(_02024_, _01905_, _01827_);
    xnor _08712_(_02025_, _01889_, _01828_);
    or _08713_(_02026_, _02025_, _01908_);
    and _08714_(_02027_, _02026_, _02024_);
    nand _08715_(_02029_, _02027_, modulus[4]);
    or _08716_(_02030_, _02029_, _02023_);
    and _08717_(_02031_, _02030_, _02022_);
    nor _08718_(_02032_, _02031_, _02014_);
    not _08719_(_02033_, _02032_);
    nand _08720_(_02034_, _02033_, _02012_);
    xor _08721_(_02035_, _02027_, _00429_);
    or _08722_(_02036_, _02035_, _02023_);
    or _08723_(_02037_, _02036_, _02014_);
    or _08724_(_02038_, _01905_, _01837_);
    or _08725_(_02040_, _01843_, modulus[0]);
    nand _08726_(_02041_, _02040_, _01884_);
    xor _08727_(_02042_, _02041_, _01838_);
    or _08728_(_02043_, _02042_, _01908_);
    and _08729_(_02044_, _02043_, _02038_);
    nand _08730_(_02045_, _02044_, modulus[3]);
    xor _08731_(_02046_, _02044_, _00309_);
    or _08732_(_02047_, _01905_, _01842_);
    xor _08733_(_02048_, _01843_, _05927_);
    or _08734_(_02049_, _02048_, _01908_);
    and _08735_(_02051_, _02049_, _02047_);
    nand _08736_(_02052_, _02051_, modulus[2]);
    or _08737_(_02053_, _02052_, _02046_);
    and _08738_(_02054_, _02053_, _02045_);
    xor _08739_(_02055_, _02051_, _00183_);
    or _08740_(_02056_, _02055_, _02046_);
    and _08741_(_02057_, _01905_, modulus[0]);
    or _08742_(_02058_, _02057_, _06035_);
    xor _08743_(_02059_, _02057_, modulus[1]);
    and _08744_(_02060_, _05927_, base[0]);
    or _08745_(_02062_, _02060_, _02059_);
    and _08746_(_02063_, _02062_, _02058_);
    or _08747_(_02064_, _02063_, _02056_);
    and _08748_(_02065_, _02064_, _02054_);
    nor _08749_(_02066_, _02065_, _02037_);
    or _08750_(_02067_, _02066_, _02034_);
    nand _08751_(_02068_, _02067_, _01993_);
    nand _08752_(_02069_, _02068_, _01988_);
    not _08753_(_02070_, _02037_);
    xor _08754_(_02071_, modulus[0], base[0]);
    nor _08755_(_02073_, _02071_, _02059_);
    not _08756_(_02074_, _02073_);
    nor _08757_(_02075_, _02074_, _02056_);
    and _08758_(_02076_, _02075_, _02070_);
    and _08759_(_02077_, _02076_, _01993_);
    not _08760_(_02078_, _02077_);
    and _08761_(_02079_, _02078_, _02069_);
    nor _08762_(_02080_, exp_counter[3], exp_counter[2]);
    nor _08763_(_02081_, exp_counter[1], exp_counter[0]);
    and _08764_(_02082_, _02081_, _02080_);
    not _08765_(_02084_, _02082_);
    and _08766_(_02085_, _02084_, _02079_);
    and _08767_(_02086_, _02085_, _01171_);
    nor _08768_(_02087_, rsa_start, rsa_active);
    and _08769_(_02088_, _02082_, _01171_);
    nor _08770_(_02089_, _02088_, _02087_);
    not _08771_(_02090_, _02089_);
    nor _08772_(_02091_, _02090_, _02086_);
    nor _08773_(_02092_, _02091_, _01138_);
    not _08774_(_02093_, _01160_);
    not _08775_(_02095_, _02079_);
    and _08776_(_02096_, _02095_, _02071_);
    and _08777_(_02097_, _02096_, _02084_);
    and _08778_(_02098_, _02097_, rsa_active);
    and _08779_(_02099_, _02098_, _02093_);
    and _08780_(_02100_, _01160_, message[0]);
    or _08781_(_02101_, _02100_, _02099_);
    and _08782_(_02102_, _02101_, _02091_);
    or _08783_(_00055_, _02102_, _02092_);
    and _08784_(_02103_, _02084_, _01171_);
    and _08785_(_02105_, _02103_, rsa_done);
    and _08786_(_02106_, _02082_, rsa_active);
    and _08787_(_02107_, _02106_, _02093_);
    not _08788_(_02108_, _02107_);
    nor _08789_(_02109_, _02108_, _02103_);
    or _08790_(_00056_, _02109_, _02105_);
    not _08791_(_02110_, _02088_);
    nor _08792_(_02111_, _01149_, exp_counter[0]);
    nor _08793_(_02112_, _02082_, _01160_);
    and _08794_(_02113_, _02112_, _02111_);
    nor _08795_(_02115_, _02113_, _02087_);
    and _08796_(_02116_, _02115_, _02110_);
    not _08797_(_02117_, _02116_);
    and _08798_(_02118_, _02117_, accumulator[0]);
    and _08799_(_02119_, accumulator[0], base[0]);
    not _08800_(_02120_, _02119_);
    and _08801_(_02121_, base[3], accumulator[12]);
    and _08802_(_02122_, base[2], accumulator[13]);
    xnor _08803_(_02123_, _02122_, _02121_);
    and _08804_(_02124_, base[1], accumulator[14]);
    xor _08805_(_02126_, _02124_, _02123_);
    and _08806_(_02127_, base[3], accumulator[11]);
    and _08807_(_02128_, base[2], accumulator[12]);
    nand _08808_(_02129_, _02128_, _02127_);
    and _08809_(_02130_, base[1], accumulator[13]);
    not _08810_(_02131_, _02130_);
    xnor _08811_(_02132_, _02128_, _02127_);
    or _08812_(_02133_, _02132_, _02131_);
    and _08813_(_02134_, _02133_, _02129_);
    xnor _08814_(_02135_, _02134_, _02126_);
    nand _08815_(_02137_, accumulator[15], base[0]);
    and _08816_(_02138_, base[4], accumulator[11]);
    xor _08817_(_02139_, _02138_, _02137_);
    and _08818_(_02140_, base[5], accumulator[10]);
    xor _08819_(_02141_, _02140_, _02139_);
    xnor _08820_(_02142_, _02141_, _02135_);
    xor _08821_(_02143_, _02132_, _02130_);
    and _08822_(_02144_, base[3], accumulator[10]);
    and _08823_(_02145_, base[2], accumulator[11]);
    nand _08824_(_02146_, _02145_, _02144_);
    and _08825_(_02148_, base[1], accumulator[12]);
    not _08826_(_02149_, _02148_);
    xnor _08827_(_02150_, _02145_, _02144_);
    or _08828_(_02151_, _02150_, _02149_);
    and _08829_(_02152_, _02151_, _02146_);
    or _08830_(_02153_, _02152_, _02143_);
    and _08831_(_02154_, accumulator[14], base[0]);
    and _08832_(_02155_, base[4], accumulator[10]);
    xnor _08833_(_02156_, _02155_, _02154_);
    and _08834_(_02157_, base[5], accumulator[9]);
    xor _08835_(_02159_, _02157_, _02156_);
    xnor _08836_(_02160_, _02152_, _02143_);
    or _08837_(_02161_, _02160_, _02159_);
    and _08838_(_02162_, _02161_, _02153_);
    xnor _08839_(_02163_, _02162_, _02142_);
    nand _08840_(_02164_, _02155_, _02154_);
    not _08841_(_02165_, _02157_);
    or _08842_(_02166_, _02165_, _02156_);
    and _08843_(_02167_, _02166_, _02164_);
    nand _08844_(_02168_, base[6], accumulator[9]);
    and _08845_(_02170_, base[7], accumulator[8]);
    xor _08846_(_02171_, _02170_, _02168_);
    and _08847_(_02172_, base[8], accumulator[7]);
    xor _08848_(_02173_, _02172_, _02171_);
    xor _08849_(_02174_, _02173_, _02167_);
    and _08850_(_02175_, base[6], accumulator[8]);
    and _08851_(_02176_, base[7], accumulator[7]);
    nand _08852_(_02177_, _02176_, _02175_);
    and _08853_(_02178_, base[8], accumulator[6]);
    not _08854_(_02179_, _02178_);
    xnor _08855_(_02181_, _02176_, _02175_);
    or _08856_(_02182_, _02181_, _02179_);
    and _08857_(_02183_, _02182_, _02177_);
    xor _08858_(_02184_, _02183_, _02174_);
    xnor _08859_(_02185_, _02184_, _02163_);
    xnor _08860_(_02186_, _02160_, _02159_);
    xor _08861_(_02187_, _02150_, _02148_);
    and _08862_(_02188_, base[3], accumulator[9]);
    and _08863_(_02189_, base[2], accumulator[10]);
    nand _08864_(_02190_, _02189_, _02188_);
    and _08865_(_02192_, base[1], accumulator[11]);
    not _08866_(_02193_, _02192_);
    xnor _08867_(_02194_, _02189_, _02188_);
    or _08868_(_02195_, _02194_, _02193_);
    and _08869_(_02196_, _02195_, _02190_);
    or _08870_(_02197_, _02196_, _02187_);
    and _08871_(_02198_, accumulator[13], base[0]);
    and _08872_(_02199_, base[4], accumulator[9]);
    xnor _08873_(_02200_, _02199_, _02198_);
    and _08874_(_02201_, base[5], accumulator[8]);
    xor _08875_(_02203_, _02201_, _02200_);
    xnor _08876_(_02204_, _02196_, _02187_);
    or _08877_(_02205_, _02204_, _02203_);
    and _08878_(_02206_, _02205_, _02197_);
    or _08879_(_02207_, _02206_, _02186_);
    and _08880_(_02208_, _02199_, _02198_);
    not _08881_(_02209_, _02201_);
    nor _08882_(_02210_, _02209_, _02200_);
    nor _08883_(_02211_, _02210_, _02208_);
    xor _08884_(_02212_, _02181_, _02178_);
    xnor _08885_(_02214_, _02212_, _02211_);
    and _08886_(_02215_, base[6], accumulator[7]);
    and _08887_(_02216_, base[7], accumulator[6]);
    nand _08888_(_02217_, _02216_, _02215_);
    and _08889_(_02218_, base[8], accumulator[5]);
    not _08890_(_02219_, _02218_);
    xnor _08891_(_02220_, _02216_, _02215_);
    or _08892_(_02221_, _02220_, _02219_);
    and _08893_(_02222_, _02221_, _02217_);
    xnor _08894_(_02223_, _02222_, _02214_);
    xnor _08895_(_02225_, _02206_, _02186_);
    or _08896_(_02226_, _02225_, _02223_);
    and _08897_(_02227_, _02226_, _02207_);
    xnor _08898_(_02228_, _02227_, _02185_);
    or _08899_(_02229_, _02212_, _02211_);
    or _08900_(_02230_, _02222_, _02214_);
    and _08901_(_02231_, _02230_, _02229_);
    nand _08902_(_02232_, base[9], accumulator[6]);
    and _08903_(_02233_, base[10], accumulator[5]);
    xor _08904_(_02234_, _02233_, _02232_);
    and _08905_(_02236_, base[11], accumulator[4]);
    xor _08906_(_02237_, _02236_, _02234_);
    and _08907_(_02238_, base[9], accumulator[5]);
    and _08908_(_02239_, base[10], accumulator[4]);
    nand _08909_(_02240_, _02239_, _02238_);
    and _08910_(_02241_, base[11], accumulator[3]);
    not _08911_(_02242_, _02241_);
    xnor _08912_(_02243_, _02239_, _02238_);
    or _08913_(_02244_, _02243_, _02242_);
    and _08914_(_02245_, _02244_, _02240_);
    xor _08915_(_02247_, _02245_, _02237_);
    nand _08916_(_02248_, base[12], accumulator[3]);
    and _08917_(_02249_, base[13], accumulator[2]);
    xor _08918_(_02250_, _02249_, _02248_);
    and _08919_(_02251_, base[14], accumulator[1]);
    xor _08920_(_02252_, _02251_, _02250_);
    xor _08921_(_02253_, _02252_, _02247_);
    xor _08922_(_02254_, _02253_, _02231_);
    xor _08923_(_02255_, _02243_, _02241_);
    and _08924_(_02256_, base[9], accumulator[4]);
    and _08925_(_02258_, base[10], accumulator[3]);
    nand _08926_(_02259_, _02258_, _02256_);
    and _08927_(_02260_, base[11], accumulator[2]);
    not _08928_(_02261_, _02260_);
    xnor _08929_(_02262_, _02258_, _02256_);
    or _08930_(_02263_, _02262_, _02261_);
    and _08931_(_02264_, _02263_, _02259_);
    or _08932_(_02265_, _02264_, _02255_);
    and _08933_(_02266_, base[12], accumulator[2]);
    and _08934_(_02267_, base[13], accumulator[1]);
    xnor _08935_(_02269_, _02267_, _02266_);
    and _08936_(_02270_, base[14], accumulator[0]);
    xor _08937_(_02271_, _02270_, _02269_);
    xnor _08938_(_02272_, _02264_, _02255_);
    or _08939_(_02273_, _02272_, _02271_);
    and _08940_(_02274_, _02273_, _02265_);
    xor _08941_(_02275_, _02274_, _02254_);
    xnor _08942_(_02276_, _02275_, _02228_);
    xnor _08943_(_02277_, _02225_, _02223_);
    xnor _08944_(_02278_, _02204_, _02203_);
    xor _08945_(_02280_, _02194_, _02192_);
    and _08946_(_02281_, base[3], accumulator[8]);
    and _08947_(_02282_, base[2], accumulator[9]);
    nand _08948_(_02283_, _02282_, _02281_);
    and _08949_(_02284_, base[1], accumulator[10]);
    not _08950_(_02285_, _02284_);
    xnor _08951_(_02286_, _02282_, _02281_);
    or _08952_(_02287_, _02286_, _02285_);
    and _08953_(_02288_, _02287_, _02283_);
    or _08954_(_02289_, _02288_, _02280_);
    and _08955_(_02291_, accumulator[12], base[0]);
    and _08956_(_02292_, base[4], accumulator[8]);
    xnor _08957_(_02293_, _02292_, _02291_);
    and _08958_(_02294_, base[5], accumulator[7]);
    xor _08959_(_02295_, _02294_, _02293_);
    xnor _08960_(_02296_, _02288_, _02280_);
    or _08961_(_02297_, _02296_, _02295_);
    and _08962_(_02298_, _02297_, _02289_);
    or _08963_(_02299_, _02298_, _02278_);
    and _08964_(_02300_, _02292_, _02291_);
    not _08965_(_02302_, _02294_);
    nor _08966_(_02303_, _02302_, _02293_);
    nor _08967_(_02304_, _02303_, _02300_);
    xor _08968_(_02305_, _02220_, _02218_);
    xnor _08969_(_02306_, _02305_, _02304_);
    and _08970_(_02307_, base[6], accumulator[6]);
    and _08971_(_02308_, base[7], accumulator[5]);
    and _08972_(_02309_, _02308_, _02307_);
    and _08973_(_02310_, base[8], accumulator[4]);
    not _08974_(_02311_, _02310_);
    xnor _08975_(_02313_, _02308_, _02307_);
    nor _08976_(_02314_, _02313_, _02311_);
    nor _08977_(_02315_, _02314_, _02309_);
    xnor _08978_(_02316_, _02315_, _02306_);
    xnor _08979_(_02317_, _02298_, _02278_);
    or _08980_(_02318_, _02317_, _02316_);
    and _08981_(_02319_, _02318_, _02299_);
    or _08982_(_02320_, _02319_, _02277_);
    nor _08983_(_02321_, _02305_, _02304_);
    nor _08984_(_02322_, _02315_, _02306_);
    nor _08985_(_02324_, _02322_, _02321_);
    xnor _08986_(_02325_, _02272_, _02271_);
    xnor _08987_(_02326_, _02325_, _02324_);
    xor _08988_(_02327_, _02262_, _02260_);
    and _08989_(_02328_, base[9], accumulator[3]);
    and _08990_(_02329_, base[10], accumulator[2]);
    and _08991_(_02330_, _02329_, _02328_);
    and _08992_(_02331_, base[11], accumulator[1]);
    not _08993_(_02332_, _02331_);
    xnor _08994_(_02333_, _02329_, _02328_);
    nor _08995_(_02335_, _02333_, _02332_);
    nor _08996_(_02336_, _02335_, _02330_);
    nor _08997_(_02337_, _02336_, _02327_);
    and _08998_(_02338_, base[12], accumulator[1]);
    and _08999_(_02339_, base[13], accumulator[0]);
    xnor _09000_(_02340_, _02339_, _02338_);
    xnor _09001_(_02341_, _02336_, _02327_);
    nor _09002_(_02342_, _02341_, _02340_);
    nor _09003_(_02343_, _02342_, _02337_);
    xnor _09004_(_02344_, _02343_, _02326_);
    xnor _09005_(_02346_, _02319_, _02277_);
    or _09006_(_02347_, _02346_, _02344_);
    and _09007_(_02348_, _02347_, _02320_);
    xnor _09008_(_02349_, _02348_, _02276_);
    nor _09009_(_02350_, _02325_, _02324_);
    nor _09010_(_02351_, _02343_, _02326_);
    or _09011_(_02352_, _02351_, _02350_);
    nand _09012_(_02353_, _02267_, _02266_);
    not _09013_(_02354_, _02270_);
    or _09014_(_02355_, _02354_, _02269_);
    and _09015_(_02357_, _02355_, _02353_);
    xor _09016_(_02358_, _02357_, _02352_);
    and _09017_(_02359_, base[15], accumulator[0]);
    xor _09018_(_02360_, _02359_, _02358_);
    xnor _09019_(_02361_, _02360_, _02349_);
    xnor _09020_(_02362_, _02346_, _02344_);
    xnor _09021_(_02363_, _02317_, _02316_);
    xnor _09022_(_02364_, _02296_, _02295_);
    xor _09023_(_02365_, _02286_, _02284_);
    and _09024_(_02366_, base[3], accumulator[7]);
    and _09025_(_02368_, base[2], accumulator[8]);
    nand _09026_(_02369_, _02368_, _02366_);
    and _09027_(_02370_, base[1], accumulator[9]);
    not _09028_(_02371_, _02370_);
    xnor _09029_(_02372_, _02368_, _02366_);
    or _09030_(_02373_, _02372_, _02371_);
    and _09031_(_02374_, _02373_, _02369_);
    or _09032_(_02375_, _02374_, _02365_);
    and _09033_(_02376_, accumulator[11], base[0]);
    and _09034_(_02377_, base[4], accumulator[7]);
    xnor _09035_(_02379_, _02377_, _02376_);
    and _09036_(_02380_, base[5], accumulator[6]);
    xor _09037_(_02381_, _02380_, _02379_);
    xnor _09038_(_02382_, _02374_, _02365_);
    or _09039_(_02383_, _02382_, _02381_);
    and _09040_(_02384_, _02383_, _02375_);
    or _09041_(_02385_, _02384_, _02364_);
    and _09042_(_02386_, _02377_, _02376_);
    not _09043_(_02387_, _02380_);
    nor _09044_(_02388_, _02387_, _02379_);
    nor _09045_(_02390_, _02388_, _02386_);
    xor _09046_(_02391_, _02313_, _02310_);
    xnor _09047_(_02392_, _02391_, _02390_);
    and _09048_(_02393_, base[6], accumulator[5]);
    and _09049_(_02394_, base[7], accumulator[4]);
    and _09050_(_02395_, _02394_, _02393_);
    and _09051_(_02396_, base[8], accumulator[3]);
    not _09052_(_02397_, _02396_);
    xnor _09053_(_02398_, _02394_, _02393_);
    nor _09054_(_02399_, _02398_, _02397_);
    nor _09055_(_02401_, _02399_, _02395_);
    xnor _09056_(_02402_, _02401_, _02392_);
    xnor _09057_(_02403_, _02384_, _02364_);
    or _09058_(_02404_, _02403_, _02402_);
    and _09059_(_02405_, _02404_, _02385_);
    or _09060_(_02406_, _02405_, _02363_);
    nor _09061_(_02407_, _02391_, _02390_);
    nor _09062_(_02408_, _02401_, _02392_);
    nor _09063_(_02409_, _02408_, _02407_);
    xnor _09064_(_02410_, _02341_, _02340_);
    xnor _09065_(_02412_, _02410_, _02409_);
    xor _09066_(_02413_, _02333_, _02331_);
    and _09067_(_02414_, base[9], accumulator[2]);
    and _09068_(_02415_, base[10], accumulator[1]);
    and _09069_(_02416_, _02415_, _02414_);
    and _09070_(_02417_, base[11], accumulator[0]);
    not _09071_(_02418_, _02417_);
    xnor _09072_(_02419_, _02415_, _02414_);
    nor _09073_(_02420_, _02419_, _02418_);
    nor _09074_(_02421_, _02420_, _02416_);
    nor _09075_(_02423_, _02421_, _02413_);
    and _09076_(_02424_, base[12], accumulator[0]);
    not _09077_(_02425_, _02424_);
    xnor _09078_(_02426_, _02421_, _02413_);
    nor _09079_(_02427_, _02426_, _02425_);
    nor _09080_(_02428_, _02427_, _02423_);
    xnor _09081_(_02429_, _02428_, _02412_);
    xnor _09082_(_02430_, _02405_, _02363_);
    or _09083_(_02431_, _02430_, _02429_);
    and _09084_(_02432_, _02431_, _02406_);
    or _09085_(_02434_, _02432_, _02362_);
    nor _09086_(_02435_, _02410_, _02409_);
    nor _09087_(_02436_, _02428_, _02412_);
    nor _09088_(_02437_, _02436_, _02435_);
    and _09089_(_02438_, _02339_, _02338_);
    xor _09090_(_02439_, _02438_, _02437_);
    xnor _09091_(_02440_, _02432_, _02362_);
    or _09092_(_02441_, _02440_, _02439_);
    and _09093_(_02442_, _02441_, _02434_);
    xnor _09094_(_02443_, _02442_, _02361_);
    not _09095_(_02445_, _02438_);
    nor _09096_(_02446_, _02445_, _02437_);
    xor _09097_(_02447_, _02446_, _02443_);
    xnor _09098_(_02448_, _02440_, _02439_);
    xnor _09099_(_02449_, _02430_, _02429_);
    xnor _09100_(_02450_, _02403_, _02402_);
    xor _09101_(_02451_, _02382_, _02381_);
    not _09102_(_02452_, _02451_);
    xor _09103_(_02453_, _02372_, _02371_);
    not _09104_(_02454_, _02453_);
    nand _09105_(_02456_, base[3], accumulator[6]);
    nand _09106_(_02457_, base[2], accumulator[7]);
    or _09107_(_02458_, _02457_, _02456_);
    nand _09108_(_02459_, base[1], accumulator[8]);
    xnor _09109_(_02460_, _02457_, _02456_);
    or _09110_(_02461_, _02460_, _02459_);
    and _09111_(_02462_, _02461_, _02458_);
    or _09112_(_02463_, _02462_, _02454_);
    and _09113_(_02464_, accumulator[10], base[0]);
    and _09114_(_02465_, base[4], accumulator[6]);
    xnor _09115_(_02467_, _02465_, _02464_);
    and _09116_(_02468_, base[5], accumulator[5]);
    xor _09117_(_02469_, _02468_, _02467_);
    xor _09118_(_02470_, _02462_, _02453_);
    or _09119_(_02471_, _02470_, _02469_);
    and _09120_(_02472_, _02471_, _02463_);
    nor _09121_(_02473_, _02472_, _02452_);
    not _09122_(_02474_, _02473_);
    and _09123_(_02475_, _02465_, _02464_);
    not _09124_(_02476_, _02475_);
    not _09125_(_02478_, _02468_);
    or _09126_(_02479_, _02478_, _02467_);
    and _09127_(_02480_, _02479_, _02476_);
    xor _09128_(_02481_, _02398_, _02396_);
    xor _09129_(_02482_, _02481_, _02480_);
    and _09130_(_02483_, base[6], accumulator[4]);
    and _09131_(_02484_, base[7], accumulator[3]);
    and _09132_(_02485_, _02484_, _02483_);
    and _09133_(_02486_, base[8], accumulator[2]);
    not _09134_(_02487_, _02486_);
    xnor _09135_(_02489_, _02484_, _02483_);
    nor _09136_(_02490_, _02489_, _02487_);
    nor _09137_(_02491_, _02490_, _02485_);
    xor _09138_(_02492_, _02491_, _02482_);
    xor _09139_(_02493_, _02472_, _02451_);
    or _09140_(_02494_, _02493_, _02492_);
    and _09141_(_02495_, _02494_, _02474_);
    nor _09142_(_02496_, _02495_, _02450_);
    not _09143_(_02497_, _02496_);
    nor _09144_(_02498_, _02481_, _02480_);
    not _09145_(_02500_, _02491_);
    and _09146_(_02501_, _02500_, _02482_);
    nor _09147_(_02502_, _02501_, _02498_);
    xor _09148_(_02503_, _02426_, _02424_);
    not _09149_(_02504_, _02503_);
    xor _09150_(_02505_, _02504_, _02502_);
    xor _09151_(_02506_, _02419_, _02417_);
    and _09152_(_02507_, base[9], accumulator[1]);
    and _09153_(_02508_, base[10], accumulator[0]);
    and _09154_(_02509_, _02508_, _02507_);
    not _09155_(_02511_, _02509_);
    nor _09156_(_02512_, _02511_, _02506_);
    xor _09157_(_02513_, _02512_, _02505_);
    xnor _09158_(_02514_, _02495_, _02450_);
    or _09159_(_02515_, _02514_, _02513_);
    and _09160_(_02516_, _02515_, _02497_);
    nor _09161_(_02517_, _02516_, _02449_);
    nor _09162_(_02518_, _02503_, _02502_);
    not _09163_(_02519_, _02512_);
    nor _09164_(_02520_, _02519_, _02505_);
    nor _09165_(_02522_, _02520_, _02518_);
    xnor _09166_(_02523_, _02516_, _02449_);
    nor _09167_(_02524_, _02523_, _02522_);
    nor _09168_(_02525_, _02524_, _02517_);
    nor _09169_(_02526_, _02525_, _02448_);
    xor _09170_(_02527_, _02526_, _02447_);
    xnor _09171_(_02528_, _02525_, _02448_);
    not _09172_(_02529_, _02528_);
    xor _09173_(_02530_, _02523_, _02522_);
    not _09174_(_02531_, _02530_);
    xor _09175_(_02533_, _02514_, _02513_);
    not _09176_(_02534_, _02533_);
    xor _09177_(_02535_, _02493_, _02492_);
    not _09178_(_02536_, _02535_);
    xnor _09179_(_02537_, _02470_, _02469_);
    xnor _09180_(_02538_, _02460_, _02459_);
    nand _09181_(_02539_, base[3], accumulator[5]);
    nand _09182_(_02540_, base[2], accumulator[6]);
    or _09183_(_02541_, _02540_, _02539_);
    nand _09184_(_02542_, base[1], accumulator[7]);
    xnor _09185_(_02544_, _02540_, _02539_);
    or _09186_(_02545_, _02544_, _02542_);
    and _09187_(_02546_, _02545_, _02541_);
    or _09188_(_02547_, _02546_, _02538_);
    nand _09189_(_02548_, accumulator[9], base[0]);
    and _09190_(_02549_, base[4], accumulator[5]);
    xor _09191_(_02550_, _02549_, _02548_);
    and _09192_(_02551_, base[5], accumulator[4]);
    xor _09193_(_02552_, _02551_, _02550_);
    xnor _09194_(_02553_, _02546_, _02538_);
    or _09195_(_02555_, _02553_, _02552_);
    and _09196_(_02556_, _02555_, _02547_);
    or _09197_(_02557_, _02556_, _02537_);
    not _09198_(_02558_, _02548_);
    nand _09199_(_02559_, _02549_, _02558_);
    not _09200_(_02560_, _02551_);
    or _09201_(_02561_, _02560_, _02550_);
    and _09202_(_02562_, _02561_, _02559_);
    xor _09203_(_02563_, _02489_, _02486_);
    xnor _09204_(_02564_, _02563_, _02562_);
    nand _09205_(_02566_, base[6], accumulator[3]);
    not _09206_(_02567_, _02566_);
    and _09207_(_02568_, base[7], accumulator[2]);
    and _09208_(_02569_, _02568_, _02567_);
    and _09209_(_02570_, base[8], accumulator[1]);
    not _09210_(_02571_, _02570_);
    xor _09211_(_02572_, _02568_, _02566_);
    nor _09212_(_02573_, _02572_, _02571_);
    nor _09213_(_02574_, _02573_, _02569_);
    xnor _09214_(_02575_, _02574_, _02564_);
    xnor _09215_(_02577_, _02556_, _02537_);
    or _09216_(_02578_, _02577_, _02575_);
    and _09217_(_02579_, _02578_, _02557_);
    or _09218_(_02580_, _02579_, _02536_);
    nor _09219_(_02581_, _02563_, _02562_);
    nor _09220_(_02582_, _02574_, _02564_);
    or _09221_(_02583_, _02582_, _02581_);
    xor _09222_(_02584_, _02509_, _02506_);
    xor _09223_(_02585_, _02584_, _02583_);
    xor _09224_(_02586_, _02579_, _02535_);
    or _09225_(_02588_, _02586_, _02585_);
    and _09226_(_02589_, _02588_, _02580_);
    or _09227_(_02590_, _02589_, _02534_);
    not _09228_(_02591_, _02584_);
    and _09229_(_02592_, _02591_, _02583_);
    not _09230_(_02593_, _02592_);
    xor _09231_(_02594_, _02589_, _02533_);
    or _09232_(_02595_, _02594_, _02593_);
    and _09233_(_02596_, _02595_, _02590_);
    nor _09234_(_02597_, _02596_, _02531_);
    nand _09235_(_02599_, _02597_, _02529_);
    xor _09236_(_02600_, _02597_, _02528_);
    xor _09237_(_02601_, _02596_, _02530_);
    xor _09238_(_02602_, _02594_, _02593_);
    not _09239_(_02603_, _02602_);
    xnor _09240_(_02604_, _02586_, _02585_);
    xnor _09241_(_02605_, _02577_, _02575_);
    xnor _09242_(_02606_, _02553_, _02552_);
    xnor _09243_(_02607_, _02544_, _02542_);
    nand _09244_(_02608_, base[3], accumulator[4]);
    nand _09245_(_02610_, base[2], accumulator[5]);
    or _09246_(_02611_, _02610_, _02608_);
    nand _09247_(_02612_, base[1], accumulator[6]);
    xnor _09248_(_02613_, _02610_, _02608_);
    or _09249_(_02614_, _02613_, _02612_);
    and _09250_(_02615_, _02614_, _02611_);
    or _09251_(_02616_, _02615_, _02607_);
    and _09252_(_02617_, accumulator[8], base[0]);
    and _09253_(_02618_, base[4], accumulator[4]);
    xnor _09254_(_02619_, _02618_, _02617_);
    and _09255_(_02621_, base[5], accumulator[3]);
    xor _09256_(_02622_, _02621_, _02619_);
    xnor _09257_(_02623_, _02615_, _02607_);
    or _09258_(_02624_, _02623_, _02622_);
    and _09259_(_02625_, _02624_, _02616_);
    or _09260_(_02626_, _02625_, _02606_);
    nand _09261_(_02627_, _02618_, _02617_);
    nand _09262_(_02628_, base[5], accumulator[3]);
    or _09263_(_02629_, _02628_, _02619_);
    and _09264_(_02630_, _02629_, _02627_);
    xor _09265_(_02632_, _02572_, _02570_);
    xnor _09266_(_02633_, _02632_, _02630_);
    nand _09267_(_02634_, base[6], accumulator[2]);
    not _09268_(_02635_, _02634_);
    and _09269_(_02636_, base[7], accumulator[1]);
    nand _09270_(_02637_, _02636_, _02635_);
    and _09271_(_02638_, base[8], accumulator[0]);
    not _09272_(_02639_, _02638_);
    xor _09273_(_02640_, _02636_, _02634_);
    or _09274_(_02641_, _02640_, _02639_);
    and _09275_(_02643_, _02641_, _02637_);
    xnor _09276_(_02644_, _02643_, _02633_);
    xnor _09277_(_02645_, _02625_, _02606_);
    or _09278_(_02646_, _02645_, _02644_);
    and _09279_(_02647_, _02646_, _02626_);
    or _09280_(_02648_, _02647_, _02605_);
    nor _09281_(_02649_, _02632_, _02630_);
    nor _09282_(_02650_, _02643_, _02633_);
    or _09283_(_02651_, _02650_, _02649_);
    xnor _09284_(_02652_, _02508_, _02507_);
    xor _09285_(_02654_, _02652_, _02651_);
    xnor _09286_(_02655_, _02647_, _02605_);
    or _09287_(_02656_, _02655_, _02654_);
    and _09288_(_02657_, _02656_, _02648_);
    or _09289_(_02658_, _02657_, _02604_);
    not _09290_(_02659_, _02652_);
    and _09291_(_02660_, _02659_, _02651_);
    not _09292_(_02661_, _02660_);
    xnor _09293_(_02662_, _02657_, _02604_);
    or _09294_(_02663_, _02662_, _02661_);
    and _09295_(_02665_, _02663_, _02658_);
    or _09296_(_02666_, _02665_, _02603_);
    or _09297_(_02667_, _02666_, _02601_);
    xnor _09298_(_02668_, _02666_, _02601_);
    xor _09299_(_02669_, _02665_, _02602_);
    xor _09300_(_02670_, _02662_, _02660_);
    xnor _09301_(_02671_, _02655_, _02654_);
    xnor _09302_(_02672_, _02645_, _02644_);
    xnor _09303_(_02673_, _02623_, _02622_);
    xnor _09304_(_02674_, _02613_, _02612_);
    nand _09305_(_02676_, base[3], accumulator[3]);
    nand _09306_(_02677_, base[2], accumulator[4]);
    or _09307_(_02678_, _02677_, _02676_);
    nand _09308_(_02679_, base[1], accumulator[5]);
    xnor _09309_(_02680_, _02677_, _02676_);
    or _09310_(_02681_, _02680_, _02679_);
    and _09311_(_02682_, _02681_, _02678_);
    or _09312_(_02683_, _02682_, _02674_);
    and _09313_(_02684_, accumulator[7], base[0]);
    and _09314_(_02685_, base[4], accumulator[3]);
    xnor _09315_(_02687_, _02685_, _02684_);
    and _09316_(_02688_, base[5], accumulator[2]);
    xor _09317_(_02689_, _02688_, _02687_);
    xnor _09318_(_02690_, _02682_, _02674_);
    or _09319_(_02691_, _02690_, _02689_);
    and _09320_(_02692_, _02691_, _02683_);
    or _09321_(_02693_, _02692_, _02673_);
    and _09322_(_02694_, _02685_, _02684_);
    not _09323_(_02695_, _02688_);
    nor _09324_(_02696_, _02695_, _02687_);
    or _09325_(_02698_, _02696_, _02694_);
    xor _09326_(_02699_, _02640_, _02638_);
    xor _09327_(_02700_, _02699_, _02698_);
    and _09328_(_02701_, base[6], accumulator[1]);
    and _09329_(_02702_, base[7], accumulator[0]);
    and _09330_(_02703_, _02702_, _02701_);
    xor _09331_(_02704_, _02703_, _02700_);
    xnor _09332_(_02705_, _02692_, _02673_);
    or _09333_(_02706_, _02705_, _02704_);
    and _09334_(_02707_, _02706_, _02693_);
    or _09335_(_02709_, _02707_, _02672_);
    not _09336_(_02710_, _02699_);
    nand _09337_(_02711_, _02710_, _02698_);
    not _09338_(_02712_, _02703_);
    or _09339_(_02713_, _02712_, _02700_);
    and _09340_(_02714_, _02713_, _02711_);
    and _09341_(_02715_, base[9], accumulator[0]);
    xor _09342_(_02716_, _02715_, _02714_);
    xnor _09343_(_02717_, _02707_, _02672_);
    or _09344_(_02718_, _02717_, _02716_);
    and _09345_(_02720_, _02718_, _02709_);
    or _09346_(_02721_, _02720_, _02671_);
    not _09347_(_02722_, _02715_);
    or _09348_(_02723_, _02722_, _02714_);
    xnor _09349_(_02724_, _02720_, _02671_);
    or _09350_(_02725_, _02724_, _02723_);
    and _09351_(_02726_, _02725_, _02721_);
    or _09352_(_02727_, _02726_, _02670_);
    or _09353_(_02728_, _02727_, _02669_);
    or _09354_(_02729_, _02728_, _02668_);
    and _09355_(_02731_, _02729_, _02667_);
    xnor _09356_(_02732_, _02727_, _02669_);
    or _09357_(_02733_, _02732_, _02668_);
    xnor _09358_(_02734_, _02726_, _02670_);
    xor _09359_(_02735_, _02724_, _02723_);
    xnor _09360_(_02736_, _02717_, _02716_);
    xnor _09361_(_02737_, _02705_, _02704_);
    xnor _09362_(_02738_, _02690_, _02689_);
    xnor _09363_(_02739_, _02680_, _02679_);
    nand _09364_(_02740_, base[3], accumulator[2]);
    nand _09365_(_02742_, base[2], accumulator[3]);
    or _09366_(_02743_, _02742_, _02740_);
    nand _09367_(_02744_, base[1], accumulator[4]);
    xnor _09368_(_02745_, _02742_, _02740_);
    or _09369_(_02746_, _02745_, _02744_);
    and _09370_(_02747_, _02746_, _02743_);
    or _09371_(_02748_, _02747_, _02739_);
    and _09372_(_02749_, accumulator[6], base[0]);
    and _09373_(_02750_, base[4], accumulator[2]);
    xnor _09374_(_02751_, _02750_, _02749_);
    and _09375_(_02753_, base[5], accumulator[1]);
    xor _09376_(_02754_, _02753_, _02751_);
    xnor _09377_(_02755_, _02747_, _02739_);
    or _09378_(_02756_, _02755_, _02754_);
    and _09379_(_02757_, _02756_, _02748_);
    or _09380_(_02758_, _02757_, _02738_);
    and _09381_(_02759_, _02750_, _02749_);
    not _09382_(_02760_, _02753_);
    nor _09383_(_02761_, _02760_, _02751_);
    or _09384_(_02762_, _02761_, _02759_);
    xnor _09385_(_02764_, _02702_, _02701_);
    xor _09386_(_02765_, _02764_, _02762_);
    xnor _09387_(_02766_, _02757_, _02738_);
    or _09388_(_02767_, _02766_, _02765_);
    and _09389_(_02768_, _02767_, _02758_);
    or _09390_(_02769_, _02768_, _02737_);
    not _09391_(_02770_, _02764_);
    and _09392_(_02771_, _02770_, _02762_);
    not _09393_(_02772_, _02771_);
    xnor _09394_(_02773_, _02768_, _02737_);
    or _09395_(_02775_, _02773_, _02772_);
    and _09396_(_02776_, _02775_, _02769_);
    nor _09397_(_02777_, _02776_, _02736_);
    nand _09398_(_02778_, _02777_, _02735_);
    or _09399_(_02779_, _02778_, _02734_);
    xnor _09400_(_02780_, _02778_, _02734_);
    xnor _09401_(_02781_, _02777_, _02735_);
    xor _09402_(_02782_, _02776_, _02736_);
    xor _09403_(_02783_, _02773_, _02771_);
    xnor _09404_(_02784_, _02766_, _02765_);
    xnor _09405_(_02786_, _02755_, _02754_);
    xnor _09406_(_02787_, _02745_, _02744_);
    and _09407_(_02788_, base[3], accumulator[1]);
    and _09408_(_02789_, base[2], accumulator[2]);
    nand _09409_(_02790_, _02789_, _02788_);
    nand _09410_(_02791_, base[1], accumulator[3]);
    xnor _09411_(_02792_, _02789_, _02788_);
    or _09412_(_02793_, _02792_, _02791_);
    and _09413_(_02794_, _02793_, _02790_);
    or _09414_(_02795_, _02794_, _02787_);
    nand _09415_(_02797_, accumulator[5], base[0]);
    and _09416_(_02798_, base[4], accumulator[1]);
    xor _09417_(_02799_, _02798_, _02797_);
    and _09418_(_02800_, base[5], accumulator[0]);
    xor _09419_(_02801_, _02800_, _02799_);
    xnor _09420_(_02802_, _02794_, _02787_);
    or _09421_(_02803_, _02802_, _02801_);
    and _09422_(_02804_, _02803_, _02795_);
    or _09423_(_02805_, _02804_, _02786_);
    not _09424_(_02806_, _02797_);
    nand _09425_(_02808_, _02798_, _02806_);
    not _09426_(_02809_, _02800_);
    or _09427_(_02810_, _02809_, _02799_);
    and _09428_(_02811_, _02810_, _02808_);
    and _09429_(_02812_, base[6], accumulator[0]);
    xor _09430_(_02813_, _02812_, _02811_);
    xnor _09431_(_02814_, _02804_, _02786_);
    or _09432_(_02815_, _02814_, _02813_);
    and _09433_(_02816_, _02815_, _02805_);
    or _09434_(_02817_, _02816_, _02784_);
    not _09435_(_02819_, _02812_);
    nor _09436_(_02820_, _02819_, _02811_);
    not _09437_(_02821_, _02820_);
    xnor _09438_(_02822_, _02816_, _02784_);
    or _09439_(_02823_, _02822_, _02821_);
    and _09440_(_02824_, _02823_, _02817_);
    nor _09441_(_02825_, _02824_, _02783_);
    nand _09442_(_02826_, _02825_, _02782_);
    or _09443_(_02827_, _02826_, _02781_);
    or _09444_(_02828_, _02827_, _02780_);
    and _09445_(_02830_, _02828_, _02779_);
    xnor _09446_(_02831_, _02826_, _02781_);
    or _09447_(_02832_, _02831_, _02780_);
    xnor _09448_(_02833_, _02825_, _02782_);
    xor _09449_(_02834_, _02824_, _02783_);
    xor _09450_(_02835_, _02822_, _02821_);
    xor _09451_(_02836_, _02814_, _02813_);
    not _09452_(_02837_, _02836_);
    xnor _09453_(_02838_, _02802_, _02801_);
    xor _09454_(_02839_, _02792_, _02791_);
    not _09455_(_02841_, _02839_);
    nand _09456_(_02842_, base[3], accumulator[0]);
    nand _09457_(_02843_, base[2], accumulator[1]);
    or _09458_(_02844_, _02843_, _02842_);
    nand _09459_(_02845_, base[1], accumulator[2]);
    xnor _09460_(_02846_, _02843_, _02842_);
    or _09461_(_02847_, _02846_, _02845_);
    and _09462_(_02848_, _02847_, _02844_);
    or _09463_(_02849_, _02848_, _02841_);
    and _09464_(_02850_, accumulator[4], base[0]);
    and _09465_(_02852_, base[4], accumulator[0]);
    xnor _09466_(_02853_, _02852_, _02850_);
    xor _09467_(_02854_, _02848_, _02839_);
    or _09468_(_02855_, _02854_, _02853_);
    and _09469_(_02856_, _02855_, _02849_);
    or _09470_(_02857_, _02856_, _02838_);
    and _09471_(_02858_, _02852_, _02850_);
    not _09472_(_02859_, _02858_);
    xnor _09473_(_02860_, _02856_, _02838_);
    or _09474_(_02861_, _02860_, _02859_);
    and _09475_(_02863_, _02861_, _02857_);
    nor _09476_(_02864_, _02863_, _02837_);
    and _09477_(_02865_, _02864_, _02835_);
    nand _09478_(_02866_, _02865_, _02834_);
    or _09479_(_02867_, _02866_, _02833_);
    xnor _09480_(_02868_, _02866_, _02833_);
    xnor _09481_(_02869_, _02865_, _02834_);
    xor _09482_(_02870_, _02864_, _02835_);
    xor _09483_(_02871_, _02863_, _02837_);
    xor _09484_(_02872_, _02860_, _02858_);
    xnor _09485_(_02874_, _02854_, _02853_);
    xnor _09486_(_02875_, _02846_, _02845_);
    and _09487_(_02876_, base[1], accumulator[1]);
    and _09488_(_02877_, base[2], accumulator[0]);
    and _09489_(_02878_, _02877_, _02876_);
    not _09490_(_02879_, _02878_);
    nor _09491_(_02880_, _02879_, _02875_);
    and _09492_(_02881_, accumulator[3], base[0]);
    not _09493_(_02882_, _02881_);
    xor _09494_(_02883_, _02878_, _02875_);
    nor _09495_(_02885_, _02883_, _02882_);
    nor _09496_(_02886_, _02885_, _02880_);
    nor _09497_(_02887_, _02886_, _02874_);
    not _09498_(_02888_, _02887_);
    nor _09499_(_02889_, _02888_, _02872_);
    and _09500_(_02890_, _02889_, _02871_);
    nand _09501_(_02891_, _02890_, _02870_);
    or _09502_(_02892_, _02891_, _02869_);
    or _09503_(_02893_, _02892_, _02868_);
    and _09504_(_02894_, _02893_, _02867_);
    or _09505_(_02896_, _02894_, _02832_);
    and _09506_(_02897_, _02896_, _02830_);
    xnor _09507_(_02898_, _02891_, _02869_);
    or _09508_(_02899_, _02898_, _02868_);
    or _09509_(_02900_, _02899_, _02832_);
    xnor _09510_(_02901_, _02890_, _02870_);
    xor _09511_(_02902_, _02889_, _02871_);
    xor _09512_(_02903_, _02887_, _02872_);
    xnor _09513_(_02904_, _02886_, _02874_);
    xor _09514_(_02905_, _02883_, _02881_);
    and _09515_(_02907_, accumulator[2], base[0]);
    not _09516_(_02908_, _02907_);
    xnor _09517_(_02909_, _02877_, _02876_);
    nor _09518_(_02910_, _02909_, _02908_);
    not _09519_(_02911_, _02910_);
    nor _09520_(_02912_, _02911_, _02905_);
    not _09521_(_02913_, _02912_);
    nor _09522_(_02914_, _02913_, _02904_);
    not _09523_(_02915_, _02914_);
    nor _09524_(_02916_, _02915_, _02903_);
    and _09525_(_02918_, _02916_, _02902_);
    not _09526_(_02919_, _02918_);
    or _09527_(_02920_, _02919_, _02901_);
    xor _09528_(_02921_, _02918_, _02901_);
    xnor _09529_(_02922_, _02916_, _02902_);
    xor _09530_(_02923_, _02914_, _02903_);
    xor _09531_(_02924_, _02912_, _02904_);
    not _09532_(_02925_, _02924_);
    xor _09533_(_02926_, _02910_, _02905_);
    xor _09534_(_02927_, _02909_, _02907_);
    and _09535_(_02929_, accumulator[1], base[0]);
    and _09536_(_02930_, base[1], accumulator[0]);
    nand _09537_(_02931_, _02930_, _02929_);
    or _09538_(_02932_, _02931_, _02927_);
    nor _09539_(_02933_, _02932_, _02926_);
    nand _09540_(_02934_, _02933_, _02925_);
    or _09541_(_02935_, _02934_, _02923_);
    or _09542_(_02936_, _02935_, _02922_);
    or _09543_(_02937_, _02936_, _02921_);
    and _09544_(_02938_, _02937_, _02920_);
    or _09545_(_02940_, _02938_, _02900_);
    and _09546_(_02941_, _02940_, _02897_);
    or _09547_(_02942_, _02941_, _02733_);
    and _09548_(_02943_, _02942_, _02731_);
    or _09549_(_02944_, _02943_, _02600_);
    and _09550_(_02945_, _02944_, _02599_);
    xnor _09551_(_02946_, _02945_, _02527_);
    or _09552_(_02947_, _02938_, _02899_);
    and _09553_(_02948_, _02947_, _02894_);
    or _09554_(_02949_, _02948_, _02831_);
    and _09555_(_02951_, _02949_, _02827_);
    xnor _09556_(_02952_, _02951_, _02780_);
    xnor _09557_(_02953_, _02948_, _02831_);
    and _09558_(_02954_, _02953_, _02952_);
    or _09559_(_02955_, _02938_, _02898_);
    and _09560_(_02956_, _02955_, _02892_);
    xnor _09561_(_02957_, _02956_, _02868_);
    xnor _09562_(_02958_, _02938_, _02898_);
    and _09563_(_02959_, _02958_, _02957_);
    and _09564_(_02960_, _02959_, _02954_);
    not _09565_(_02962_, _02960_);
    or _09566_(_02963_, _02941_, _02732_);
    and _09567_(_02964_, _02963_, _02728_);
    xnor _09568_(_02965_, _02964_, _02668_);
    xnor _09569_(_02966_, _02941_, _02732_);
    nand _09570_(_02967_, _02966_, _02965_);
    xor _09571_(_02968_, _02946_, _05927_);
    xnor _09572_(_02969_, _02943_, _02600_);
    not _09573_(_02970_, _02969_);
    or _09574_(_02971_, _02970_, _02968_);
    or _09575_(_02973_, _02971_, _02967_);
    or _09576_(_02974_, _02973_, _02962_);
    xnor _09577_(_02975_, _02936_, _02921_);
    xnor _09578_(_02976_, _02935_, _02922_);
    and _09579_(_02977_, _02976_, _02975_);
    and _09580_(_02978_, _02933_, _02925_);
    xor _09581_(_02979_, _02978_, _02923_);
    xor _09582_(_02980_, _02933_, _02924_);
    and _09583_(_02981_, _02980_, _02979_);
    and _09584_(_02982_, _02981_, _02977_);
    xnor _09585_(_02984_, _02932_, _02926_);
    xnor _09586_(_02985_, _02931_, _02927_);
    and _09587_(_02986_, _02985_, _02984_);
    xnor _09588_(_02987_, _02930_, _02929_);
    and _09589_(_02988_, _02987_, _02120_);
    and _09590_(_02989_, _02988_, _02986_);
    and _09591_(_02990_, _02989_, _02982_);
    not _09592_(_02991_, _02990_);
    nor _09593_(_02992_, _02991_, _02974_);
    nand _09594_(_02993_, _02992_, _05960_);
    or _09595_(_02995_, _02946_, modulus[0]);
    or _09596_(_02996_, _02969_, _02968_);
    and _09597_(_02997_, _02996_, _02995_);
    and _09598_(_02998_, _02966_, _02965_);
    or _09599_(_02999_, _02998_, _02971_);
    and _09600_(_03000_, _02999_, _02997_);
    and _09601_(_03001_, _02953_, _02952_);
    and _09602_(_03002_, _02958_, _02957_);
    not _09603_(_03003_, _03002_);
    nand _09604_(_03004_, _03003_, _02954_);
    and _09605_(_03006_, _03004_, _03001_);
    or _09606_(_03007_, _03006_, _02973_);
    and _09607_(_03008_, _03007_, _03000_);
    and _09608_(_03009_, _02976_, _02975_);
    nand _09609_(_03010_, _02980_, _02979_);
    nand _09610_(_03011_, _03010_, _02977_);
    and _09611_(_03012_, _03011_, _03009_);
    nand _09612_(_03013_, _02981_, _02977_);
    and _09613_(_03014_, _03013_, _03012_);
    or _09614_(_03015_, _03014_, _02974_);
    nand _09615_(_03017_, _03015_, _03008_);
    and _09616_(_03018_, _03017_, _05952_);
    and _09617_(_03019_, _03018_, _05955_);
    and _09618_(_03020_, _03019_, _05957_);
    nand _09619_(_03021_, _03020_, _05956_);
    nand _09620_(_03022_, _03021_, _02993_);
    or _09621_(_03023_, _03022_, _02946_);
    and _09622_(_03024_, _03021_, _02993_);
    not _09623_(_03025_, _03014_);
    nand _09624_(_03026_, _03025_, _02960_);
    and _09625_(_03028_, _03026_, _03006_);
    or _09626_(_03029_, _03028_, _02967_);
    and _09627_(_03030_, _03029_, _02998_);
    nand _09628_(_03031_, _03030_, _02969_);
    xor _09629_(_03032_, _03031_, _02968_);
    or _09630_(_03033_, _03032_, _03024_);
    and _09631_(_03034_, _03033_, _03023_);
    or _09632_(_03035_, _03022_, _02952_);
    nand _09633_(_03036_, _03025_, _02959_);
    and _09634_(_03037_, _03036_, _03002_);
    and _09635_(_03039_, _03037_, _02953_);
    xor _09636_(_03040_, _03039_, _02952_);
    or _09637_(_03041_, _03040_, _03024_);
    nand _09638_(_03042_, _03041_, _03035_);
    or _09639_(_03043_, _03022_, _02953_);
    xor _09640_(_03044_, _03037_, _02953_);
    or _09641_(_03045_, _03044_, _03024_);
    nand _09642_(_03046_, _03045_, _03043_);
    or _09643_(_03047_, _03046_, _03042_);
    or _09644_(_03048_, _03022_, _02957_);
    and _09645_(_03050_, _03014_, _02958_);
    xor _09646_(_03051_, _03050_, _02957_);
    or _09647_(_03052_, _03051_, _03024_);
    and _09648_(_03053_, _03052_, _03048_);
    or _09649_(_03054_, _03022_, _02958_);
    xor _09650_(_03055_, _03014_, _02958_);
    or _09651_(_03056_, _03055_, _03024_);
    and _09652_(_03057_, _03056_, _03054_);
    nand _09653_(_03058_, _03057_, _03053_);
    or _09654_(_03059_, _03058_, _03047_);
    or _09655_(_03061_, _03022_, _02965_);
    and _09656_(_03062_, _03028_, _02966_);
    xor _09657_(_03063_, _03062_, _02965_);
    or _09658_(_03064_, _03063_, _03024_);
    nand _09659_(_03065_, _03064_, _03061_);
    or _09660_(_03066_, _03022_, _02966_);
    xor _09661_(_03067_, _03028_, _02966_);
    or _09662_(_03068_, _03067_, _03024_);
    nand _09663_(_03069_, _03068_, _03066_);
    or _09664_(_03070_, _03069_, _03065_);
    xor _09665_(_03072_, _03034_, _06035_);
    or _09666_(_03073_, _03022_, _02969_);
    xor _09667_(_03074_, _03030_, _02969_);
    or _09668_(_03075_, _03074_, _03024_);
    and _09669_(_03076_, _03075_, _03073_);
    xor _09670_(_03077_, _03076_, _05927_);
    or _09671_(_03078_, _03077_, _03072_);
    or _09672_(_03079_, _03078_, _03070_);
    or _09673_(_03080_, _03079_, _03059_);
    not _09674_(_03081_, _02989_);
    or _09675_(_03083_, _03022_, _02975_);
    and _09676_(_03084_, _02980_, _02979_);
    nor _09677_(_03085_, _03084_, _03010_);
    and _09678_(_03086_, _03085_, _02976_);
    xor _09679_(_03087_, _03086_, _02975_);
    or _09680_(_03088_, _03087_, _03024_);
    and _09681_(_03089_, _03088_, _03083_);
    or _09682_(_03090_, _03022_, _02976_);
    xor _09683_(_03091_, _03085_, _02976_);
    or _09684_(_03092_, _03091_, _03024_);
    and _09685_(_03094_, _03092_, _03090_);
    nand _09686_(_03095_, _03094_, _03089_);
    nand _09687_(_03096_, _02980_, _02979_);
    or _09688_(_03097_, _03096_, _03095_);
    or _09689_(_03098_, _03097_, _03081_);
    nor _09690_(_03099_, _03098_, _03080_);
    nand _09691_(_03100_, _03099_, _06076_);
    or _09692_(_03101_, _03034_, modulus[1]);
    or _09693_(_03102_, _03076_, modulus[0]);
    or _09694_(_03103_, _03102_, _03072_);
    and _09695_(_03105_, _03103_, _03101_);
    and _09696_(_03106_, _03064_, _03061_);
    and _09697_(_03107_, _03068_, _03066_);
    and _09698_(_03108_, _03107_, _03106_);
    or _09699_(_03109_, _03108_, _03078_);
    and _09700_(_03110_, _03109_, _03105_);
    and _09701_(_03111_, _03041_, _03035_);
    and _09702_(_03112_, _03045_, _03043_);
    and _09703_(_03113_, _03112_, _03111_);
    and _09704_(_03114_, _03057_, _03053_);
    or _09705_(_03116_, _03114_, _03047_);
    and _09706_(_03117_, _03116_, _03113_);
    or _09707_(_03118_, _03117_, _03079_);
    and _09708_(_03119_, _03118_, _03110_);
    and _09709_(_03120_, _03094_, _03089_);
    and _09710_(_03121_, _02980_, _02979_);
    or _09711_(_03122_, _03121_, _03095_);
    and _09712_(_03123_, _03122_, _03120_);
    not _09713_(_03124_, _02986_);
    and _09714_(_03125_, _02985_, _02984_);
    and _09715_(_03127_, _03125_, _03124_);
    or _09716_(_03128_, _03097_, _03127_);
    and _09717_(_03129_, _03128_, _03123_);
    or _09718_(_03130_, _03129_, _03080_);
    nand _09719_(_03131_, _03130_, _03119_);
    and _09720_(_03132_, _03131_, _06070_);
    and _09721_(_03133_, _03132_, _06074_);
    nand _09722_(_03134_, _03133_, _06071_);
    nand _09723_(_03135_, _03134_, _03100_);
    or _09724_(_03136_, _03135_, _03034_);
    and _09725_(_03138_, _03134_, _03100_);
    or _09726_(_03139_, _03129_, _03059_);
    and _09727_(_03140_, _03139_, _03117_);
    or _09728_(_03141_, _03140_, _03070_);
    and _09729_(_03142_, _03141_, _03108_);
    or _09730_(_03143_, _03142_, _03077_);
    nand _09731_(_03144_, _03143_, _03102_);
    xor _09732_(_03145_, _03144_, _03072_);
    or _09733_(_03146_, _03145_, _03138_);
    and _09734_(_03147_, _03146_, _03136_);
    or _09735_(_03149_, _03135_, _03111_);
    or _09736_(_03150_, _03129_, _03058_);
    and _09737_(_03151_, _03150_, _03114_);
    and _09738_(_03152_, _03151_, _03112_);
    xor _09739_(_03153_, _03152_, _03042_);
    nand _09740_(_03154_, _03153_, _03135_);
    nand _09741_(_03155_, _03154_, _03149_);
    or _09742_(_03156_, _03135_, _03112_);
    xor _09743_(_03157_, _03151_, _03046_);
    nand _09744_(_03158_, _03157_, _03135_);
    nand _09745_(_03160_, _03158_, _03156_);
    or _09746_(_03161_, _03160_, _03155_);
    or _09747_(_03162_, _03135_, _03053_);
    and _09748_(_03163_, _03129_, _03057_);
    xor _09749_(_03164_, _03163_, _03053_);
    or _09750_(_03165_, _03164_, _03138_);
    and _09751_(_03166_, _03165_, _03162_);
    or _09752_(_03167_, _03135_, _03057_);
    xor _09753_(_03168_, _03129_, _03057_);
    or _09754_(_03169_, _03168_, _03138_);
    and _09755_(_03171_, _03169_, _03167_);
    nand _09756_(_03172_, _03171_, _03166_);
    or _09757_(_03173_, _03172_, _03161_);
    or _09758_(_03174_, _03135_, _03106_);
    and _09759_(_03175_, _03140_, _03107_);
    xor _09760_(_03176_, _03175_, _03065_);
    nand _09761_(_03177_, _03176_, _03135_);
    and _09762_(_03178_, _03177_, _03174_);
    xor _09763_(_03179_, _03178_, _05927_);
    or _09764_(_03180_, _03135_, _03107_);
    xor _09765_(_03182_, _03140_, _03069_);
    nand _09766_(_03183_, _03182_, _03135_);
    and _09767_(_03184_, _03183_, _03180_);
    not _09768_(_03185_, _03184_);
    or _09769_(_03186_, _03185_, _03179_);
    xor _09770_(_03187_, _03147_, _00183_);
    or _09771_(_03188_, _03135_, _03076_);
    xnor _09772_(_03189_, _03142_, _03077_);
    or _09773_(_03190_, _03189_, _03138_);
    and _09774_(_03191_, _03190_, _03188_);
    xor _09775_(_03193_, _03191_, _06035_);
    or _09776_(_03194_, _03193_, _03187_);
    or _09777_(_03195_, _03194_, _03186_);
    or _09778_(_03196_, _03195_, _03173_);
    or _09779_(_03197_, _03135_, _03089_);
    nand _09780_(_03198_, _02980_, _02979_);
    and _09781_(_03199_, _03198_, _03121_);
    and _09782_(_03200_, _03199_, _03094_);
    xor _09783_(_03201_, _03200_, _03089_);
    or _09784_(_03202_, _03201_, _03138_);
    nand _09785_(_03204_, _03202_, _03197_);
    or _09786_(_03205_, _03135_, _03094_);
    xor _09787_(_03206_, _03199_, _03094_);
    or _09788_(_03207_, _03206_, _03138_);
    nand _09789_(_03208_, _03207_, _03205_);
    or _09790_(_03209_, _03208_, _03204_);
    or _09791_(_03210_, _03022_, _02979_);
    xor _09792_(_03211_, _02978_, _02923_);
    or _09793_(_03212_, _03211_, _03024_);
    and _09794_(_03213_, _03212_, _03210_);
    or _09795_(_03215_, _03135_, _03213_);
    xor _09796_(_03216_, _02933_, _02924_);
    and _09797_(_03217_, _03216_, _03127_);
    xor _09798_(_03218_, _03217_, _03213_);
    or _09799_(_03219_, _03218_, _03138_);
    and _09800_(_03220_, _03219_, _03215_);
    or _09801_(_03221_, _03135_, _03216_);
    xor _09802_(_03222_, _02933_, _02924_);
    or _09803_(_03223_, _03222_, _03138_);
    and _09804_(_03224_, _03223_, _03221_);
    nand _09805_(_03226_, _03224_, _03220_);
    or _09806_(_03227_, _03226_, _03209_);
    nor _09807_(_03228_, _03227_, _03081_);
    not _09808_(_03229_, _03228_);
    nor _09809_(_03230_, _03229_, _03196_);
    nand _09810_(_03231_, _03230_, _00231_);
    or _09811_(_03232_, _03147_, modulus[2]);
    or _09812_(_03233_, _03191_, modulus[1]);
    or _09813_(_03234_, _03233_, _03187_);
    and _09814_(_03235_, _03234_, _03232_);
    or _09815_(_03237_, _03178_, modulus[0]);
    or _09816_(_03238_, _03184_, _03179_);
    and _09817_(_03239_, _03238_, _03237_);
    or _09818_(_03240_, _03239_, _03194_);
    and _09819_(_03241_, _03240_, _03235_);
    nor _09820_(_03242_, _03160_, _03155_);
    and _09821_(_03243_, _03171_, _03166_);
    or _09822_(_03244_, _03243_, _03161_);
    and _09823_(_03245_, _03244_, _03242_);
    or _09824_(_03246_, _03245_, _03195_);
    and _09825_(_03248_, _03246_, _03241_);
    nor _09826_(_03249_, _03208_, _03204_);
    and _09827_(_03250_, _03224_, _03220_);
    or _09828_(_03251_, _03250_, _03209_);
    and _09829_(_03252_, _03251_, _03249_);
    or _09830_(_03253_, _03227_, _03127_);
    and _09831_(_03254_, _03253_, _03252_);
    or _09832_(_03255_, _03254_, _03196_);
    nand _09833_(_03256_, _03255_, _03248_);
    and _09834_(_03257_, _03256_, _00228_);
    and _09835_(_03259_, _03257_, _00229_);
    nand _09836_(_03260_, _03259_, _05956_);
    nand _09837_(_03261_, _03260_, _03231_);
    or _09838_(_03262_, _03261_, _03147_);
    and _09839_(_03263_, _03260_, _03231_);
    or _09840_(_03264_, _03254_, _03173_);
    and _09841_(_03265_, _03264_, _03245_);
    or _09842_(_03266_, _03265_, _03186_);
    and _09843_(_03267_, _03266_, _03239_);
    or _09844_(_03268_, _03267_, _03193_);
    nand _09845_(_03270_, _03268_, _03233_);
    xor _09846_(_03271_, _03270_, _03187_);
    or _09847_(_03272_, _03271_, _03263_);
    and _09848_(_03273_, _03272_, _03262_);
    nand _09849_(_03274_, _03263_, _03155_);
    not _09850_(_03275_, _03160_);
    or _09851_(_03276_, _03254_, _03172_);
    and _09852_(_03277_, _03276_, _03243_);
    and _09853_(_03278_, _03277_, _03275_);
    xor _09854_(_03279_, _03278_, _03155_);
    nand _09855_(_03281_, _03279_, _03261_);
    nand _09856_(_03282_, _03281_, _03274_);
    or _09857_(_03283_, _03261_, _03275_);
    xor _09858_(_03284_, _03277_, _03275_);
    or _09859_(_03285_, _03284_, _03263_);
    nand _09860_(_03286_, _03285_, _03283_);
    or _09861_(_03287_, _03286_, _03282_);
    or _09862_(_03288_, _03261_, _03166_);
    and _09863_(_03289_, _03254_, _03171_);
    xor _09864_(_03290_, _03289_, _03166_);
    or _09865_(_03292_, _03290_, _03263_);
    and _09866_(_03293_, _03292_, _03288_);
    or _09867_(_03294_, _03261_, _03171_);
    xor _09868_(_03295_, _03254_, _03171_);
    or _09869_(_03296_, _03295_, _03263_);
    and _09870_(_03297_, _03296_, _03294_);
    nand _09871_(_03298_, _03297_, _03293_);
    or _09872_(_03299_, _03298_, _03287_);
    or _09873_(_03300_, _03261_, _03178_);
    and _09874_(_03301_, _03265_, _03184_);
    xor _09875_(_03303_, _03301_, _03179_);
    nand _09876_(_03304_, _03303_, _03261_);
    and _09877_(_03305_, _03304_, _03300_);
    xor _09878_(_03306_, _03305_, _06035_);
    or _09879_(_03307_, _03261_, _03184_);
    xor _09880_(_03308_, _03265_, _03185_);
    nand _09881_(_03309_, _03308_, _03261_);
    and _09882_(_03310_, _03309_, _03307_);
    xor _09883_(_03311_, _03310_, _05927_);
    or _09884_(_03312_, _03311_, _03306_);
    xor _09885_(_03314_, _03273_, _00309_);
    or _09886_(_03315_, _03261_, _03191_);
    xnor _09887_(_03316_, _03267_, _03193_);
    or _09888_(_03317_, _03316_, _03263_);
    and _09889_(_03318_, _03317_, _03315_);
    xor _09890_(_03319_, _03318_, _00183_);
    or _09891_(_03320_, _03319_, _03314_);
    or _09892_(_03321_, _03320_, _03312_);
    nor _09893_(_03322_, _03321_, _03299_);
    not _09894_(_03323_, _03204_);
    or _09895_(_03325_, _03261_, _03323_);
    not _09896_(_03326_, _03208_);
    or _09897_(_03327_, _03226_, _03127_);
    and _09898_(_03328_, _03327_, _03250_);
    and _09899_(_03329_, _03328_, _03326_);
    xor _09900_(_03330_, _03329_, _03323_);
    or _09901_(_03331_, _03330_, _03263_);
    and _09902_(_03332_, _03331_, _03325_);
    or _09903_(_03333_, _03261_, _03326_);
    xor _09904_(_03334_, _03328_, _03326_);
    or _09905_(_03336_, _03334_, _03263_);
    and _09906_(_03337_, _03336_, _03333_);
    nand _09907_(_03338_, _03337_, _03332_);
    or _09908_(_03339_, _03261_, _03220_);
    and _09909_(_03340_, _03224_, _03127_);
    xor _09910_(_03341_, _03340_, _03220_);
    or _09911_(_03342_, _03341_, _03263_);
    and _09912_(_03343_, _03342_, _03339_);
    or _09913_(_03344_, _03261_, _03224_);
    xor _09914_(_03345_, _03224_, _03127_);
    or _09915_(_03347_, _03345_, _03263_);
    and _09916_(_03348_, _03347_, _03344_);
    nand _09917_(_03349_, _03348_, _03343_);
    nor _09918_(_03350_, _03349_, _03338_);
    and _09919_(_03351_, _03350_, _02989_);
    and _09920_(_03352_, _03351_, _03322_);
    nand _09921_(_03353_, _03352_, _00350_);
    or _09922_(_03354_, _03273_, modulus[3]);
    or _09923_(_03355_, _03318_, modulus[2]);
    or _09924_(_03356_, _03355_, _03314_);
    and _09925_(_03358_, _03356_, _03354_);
    or _09926_(_03359_, _03305_, modulus[1]);
    or _09927_(_03360_, _03310_, modulus[0]);
    or _09928_(_03361_, _03360_, _03306_);
    and _09929_(_03362_, _03361_, _03359_);
    or _09930_(_03363_, _03362_, _03320_);
    and _09931_(_03364_, _03363_, _03358_);
    nor _09932_(_03365_, _03286_, _03282_);
    and _09933_(_03366_, _03297_, _03293_);
    or _09934_(_03367_, _03366_, _03287_);
    and _09935_(_03369_, _03367_, _03365_);
    or _09936_(_03370_, _03369_, _03321_);
    and _09937_(_03371_, _03370_, _03364_);
    and _09938_(_03372_, _03337_, _03332_);
    and _09939_(_03373_, _03348_, _03343_);
    or _09940_(_03374_, _03373_, _03338_);
    and _09941_(_03375_, _03374_, _03372_);
    not _09942_(_03376_, _03127_);
    nand _09943_(_03377_, _03350_, _03376_);
    nand _09944_(_03378_, _03377_, _03375_);
    nand _09945_(_03380_, _03378_, _03322_);
    nand _09946_(_03381_, _03380_, _03371_);
    and _09947_(_03382_, _03381_, _00349_);
    nand _09948_(_03383_, _03382_, _00346_);
    nand _09949_(_03384_, _03383_, _03353_);
    or _09950_(_03385_, _03384_, _03273_);
    and _09951_(_03386_, _03377_, _03375_);
    or _09952_(_03387_, _03386_, _03299_);
    and _09953_(_03388_, _03387_, _03369_);
    or _09954_(_03389_, _03388_, _03312_);
    and _09955_(_03391_, _03389_, _03362_);
    or _09956_(_03392_, _03391_, _03319_);
    and _09957_(_03393_, _03392_, _03355_);
    xor _09958_(_03394_, _03393_, _03314_);
    nand _09959_(_03395_, _03394_, _03384_);
    and _09960_(_03396_, _03395_, _03385_);
    and _09961_(_03397_, _03383_, _03353_);
    nand _09962_(_03398_, _03397_, _03282_);
    not _09963_(_03399_, _03286_);
    or _09964_(_03400_, _03386_, _03298_);
    and _09965_(_03402_, _03400_, _03366_);
    and _09966_(_03403_, _03402_, _03399_);
    xor _09967_(_03404_, _03403_, _03282_);
    nand _09968_(_03405_, _03404_, _03384_);
    and _09969_(_03406_, _03405_, _03398_);
    xor _09970_(_03407_, _03406_, _05927_);
    or _09971_(_03408_, _03384_, _03399_);
    xor _09972_(_03409_, _03402_, _03286_);
    nand _09973_(_03410_, _03409_, _03384_);
    nand _09974_(_03411_, _03410_, _03408_);
    or _09975_(_03413_, _03411_, _03407_);
    or _09976_(_03414_, _03384_, _03293_);
    and _09977_(_03415_, _03386_, _03297_);
    xor _09978_(_03416_, _03415_, _03293_);
    or _09979_(_03417_, _03416_, _03397_);
    and _09980_(_03418_, _03417_, _03414_);
    or _09981_(_03419_, _03384_, _03297_);
    xor _09982_(_03420_, _03386_, _03297_);
    or _09983_(_03421_, _03420_, _03397_);
    and _09984_(_03422_, _03421_, _03419_);
    nand _09985_(_03424_, _03422_, _03418_);
    or _09986_(_03425_, _03424_, _03413_);
    or _09987_(_03426_, _03384_, _03305_);
    or _09988_(_03427_, _03388_, _03311_);
    and _09989_(_03428_, _03427_, _03360_);
    xor _09990_(_03429_, _03428_, _03306_);
    nand _09991_(_03430_, _03429_, _03384_);
    and _09992_(_03431_, _03430_, _03426_);
    xor _09993_(_03432_, _03431_, _00183_);
    or _09994_(_03433_, _03384_, _03310_);
    xor _09995_(_03435_, _03388_, _03311_);
    nand _09996_(_03436_, _03435_, _03384_);
    and _09997_(_03437_, _03436_, _03433_);
    xor _09998_(_03438_, _03437_, _06035_);
    or _09999_(_03439_, _03438_, _03432_);
    xor _10000_(_03440_, _03396_, _00429_);
    or _10001_(_03441_, _03384_, _03318_);
    xor _10002_(_03442_, _03391_, _03319_);
    nand _10003_(_03443_, _03442_, _03384_);
    and _10004_(_03444_, _03443_, _03441_);
    xor _10005_(_03446_, _03444_, _00309_);
    or _10006_(_03447_, _03446_, _03440_);
    or _10007_(_03448_, _03447_, _03439_);
    nor _10008_(_03449_, _03448_, _03425_);
    or _10009_(_03450_, _03384_, _03332_);
    or _10010_(_03451_, _03349_, _03127_);
    and _10011_(_03452_, _03451_, _03373_);
    and _10012_(_03453_, _03452_, _03337_);
    xor _10013_(_03454_, _03453_, _03332_);
    or _10014_(_03455_, _03454_, _03397_);
    nand _10015_(_03457_, _03455_, _03450_);
    or _10016_(_03458_, _03384_, _03337_);
    xor _10017_(_03459_, _03452_, _03337_);
    or _10018_(_03460_, _03459_, _03397_);
    nand _10019_(_03461_, _03460_, _03458_);
    or _10020_(_03462_, _03461_, _03457_);
    or _10021_(_03463_, _03384_, _03343_);
    and _10022_(_03464_, _03348_, _03127_);
    xor _10023_(_03465_, _03464_, _03343_);
    or _10024_(_03466_, _03465_, _03397_);
    and _10025_(_03468_, _03466_, _03463_);
    or _10026_(_03469_, _03384_, _03348_);
    xor _10027_(_03470_, _03348_, _03127_);
    or _10028_(_03471_, _03470_, _03397_);
    and _10029_(_03472_, _03471_, _03469_);
    nand _10030_(_03473_, _03472_, _03468_);
    nor _10031_(_03474_, _03473_, _03462_);
    and _10032_(_03475_, _03474_, _02989_);
    and _10033_(_03476_, _03475_, _03449_);
    nand _10034_(_03477_, _03476_, _00467_);
    or _10035_(_03479_, _03396_, modulus[4]);
    or _10036_(_03480_, _03444_, modulus[3]);
    or _10037_(_03481_, _03480_, _03440_);
    and _10038_(_03482_, _03481_, _03479_);
    or _10039_(_03483_, _03431_, modulus[2]);
    or _10040_(_03484_, _03437_, modulus[1]);
    or _10041_(_03485_, _03484_, _03432_);
    and _10042_(_03486_, _03485_, _03483_);
    or _10043_(_03487_, _03486_, _03447_);
    and _10044_(_03488_, _03487_, _03482_);
    or _10045_(_03490_, _03406_, modulus[0]);
    and _10046_(_03491_, _03410_, _03408_);
    or _10047_(_03492_, _03491_, _03407_);
    and _10048_(_03493_, _03492_, _03490_);
    and _10049_(_03494_, _03422_, _03418_);
    or _10050_(_03495_, _03494_, _03413_);
    and _10051_(_03496_, _03495_, _03493_);
    or _10052_(_03497_, _03496_, _03448_);
    and _10053_(_03498_, _03497_, _03488_);
    nor _10054_(_03499_, _03461_, _03457_);
    and _10055_(_03501_, _03472_, _03468_);
    or _10056_(_03502_, _03501_, _03462_);
    and _10057_(_03503_, _03502_, _03499_);
    nand _10058_(_03504_, _03474_, _03376_);
    nand _10059_(_03505_, _03504_, _03503_);
    nand _10060_(_03506_, _03505_, _03449_);
    nand _10061_(_03507_, _03506_, _03498_);
    and _10062_(_03508_, _03507_, _00466_);
    and _10063_(_03509_, _03508_, _05957_);
    nand _10064_(_03510_, _03509_, _05956_);
    nand _10065_(_03512_, _03510_, _03477_);
    or _10066_(_03513_, _03512_, _03396_);
    and _10067_(_03514_, _03504_, _03503_);
    or _10068_(_03515_, _03514_, _03425_);
    and _10069_(_03516_, _03515_, _03496_);
    or _10070_(_03517_, _03516_, _03439_);
    and _10071_(_03518_, _03517_, _03486_);
    or _10072_(_03519_, _03518_, _03446_);
    and _10073_(_03520_, _03519_, _03480_);
    xor _10074_(_03521_, _03520_, _03440_);
    nand _10075_(_03523_, _03521_, _03512_);
    and _10076_(_03524_, _03523_, _03513_);
    or _10077_(_03525_, _03512_, _03406_);
    or _10078_(_03526_, _03514_, _03424_);
    and _10079_(_03527_, _03526_, _03494_);
    and _10080_(_03528_, _03527_, _03491_);
    xor _10081_(_03529_, _03528_, _03407_);
    nand _10082_(_03530_, _03529_, _03512_);
    and _10083_(_03531_, _03530_, _03525_);
    xor _10084_(_03532_, _03531_, _06035_);
    or _10085_(_03534_, _03512_, _03491_);
    xor _10086_(_03535_, _03527_, _03411_);
    nand _10087_(_03536_, _03535_, _03512_);
    and _10088_(_03537_, _03536_, _03534_);
    xor _10089_(_03538_, _03537_, _05927_);
    or _10090_(_03539_, _03538_, _03532_);
    or _10091_(_03540_, _03512_, _03418_);
    and _10092_(_03541_, _03510_, _03477_);
    and _10093_(_03542_, _03514_, _03422_);
    xor _10094_(_03543_, _03542_, _03418_);
    or _10095_(_03545_, _03543_, _03541_);
    and _10096_(_03546_, _03545_, _03540_);
    or _10097_(_03547_, _03512_, _03422_);
    xor _10098_(_03548_, _03514_, _03422_);
    or _10099_(_03549_, _03548_, _03541_);
    and _10100_(_03550_, _03549_, _03547_);
    nand _10101_(_03551_, _03550_, _03546_);
    or _10102_(_03552_, _03551_, _03539_);
    or _10103_(_03553_, _03512_, _03431_);
    or _10104_(_03554_, _03516_, _03438_);
    and _10105_(_03556_, _03554_, _03484_);
    xor _10106_(_03557_, _03556_, _03432_);
    nand _10107_(_03558_, _03557_, _03512_);
    and _10108_(_03559_, _03558_, _03553_);
    xor _10109_(_03560_, _03559_, _00309_);
    or _10110_(_03561_, _03512_, _03437_);
    xor _10111_(_03562_, _03516_, _03438_);
    nand _10112_(_03563_, _03562_, _03512_);
    and _10113_(_03564_, _03563_, _03561_);
    xor _10114_(_03565_, _03564_, _00183_);
    or _10115_(_03567_, _03565_, _03560_);
    xor _10116_(_03568_, _03524_, _00550_);
    or _10117_(_03569_, _03512_, _03444_);
    xor _10118_(_03570_, _03518_, _03446_);
    nand _10119_(_03571_, _03570_, _03512_);
    and _10120_(_03572_, _03571_, _03569_);
    xor _10121_(_03573_, _03572_, _00429_);
    or _10122_(_03574_, _03573_, _03568_);
    or _10123_(_03575_, _03574_, _03567_);
    nor _10124_(_03576_, _03575_, _03552_);
    not _10125_(_03578_, _03457_);
    or _10126_(_03579_, _03512_, _03578_);
    not _10127_(_03580_, _03461_);
    or _10128_(_03581_, _03473_, _03127_);
    and _10129_(_03582_, _03581_, _03501_);
    and _10130_(_03583_, _03582_, _03580_);
    xor _10131_(_03584_, _03583_, _03578_);
    or _10132_(_03585_, _03584_, _03541_);
    nand _10133_(_03586_, _03585_, _03579_);
    or _10134_(_03587_, _03512_, _03580_);
    xor _10135_(_03589_, _03582_, _03580_);
    or _10136_(_03590_, _03589_, _03541_);
    nand _10137_(_03591_, _03590_, _03587_);
    or _10138_(_03592_, _03591_, _03586_);
    or _10139_(_03593_, _03512_, _03468_);
    and _10140_(_03594_, _03472_, _03127_);
    xor _10141_(_03595_, _03594_, _03468_);
    or _10142_(_03596_, _03595_, _03541_);
    and _10143_(_03597_, _03596_, _03593_);
    or _10144_(_03598_, _03512_, _03472_);
    xor _10145_(_03600_, _03472_, _03127_);
    or _10146_(_03601_, _03600_, _03541_);
    and _10147_(_03602_, _03601_, _03598_);
    nand _10148_(_03603_, _03602_, _03597_);
    nor _10149_(_03604_, _03603_, _03592_);
    and _10150_(_03605_, _03604_, _02989_);
    and _10151_(_03606_, _03605_, _03576_);
    nand _10152_(_03607_, _03606_, _00588_);
    or _10153_(_03608_, _03524_, modulus[5]);
    or _10154_(_03609_, _03572_, modulus[4]);
    or _10155_(_03611_, _03609_, _03568_);
    and _10156_(_03612_, _03611_, _03608_);
    or _10157_(_03613_, _03559_, modulus[3]);
    or _10158_(_03614_, _03564_, modulus[2]);
    or _10159_(_03615_, _03614_, _03560_);
    and _10160_(_03616_, _03615_, _03613_);
    or _10161_(_03617_, _03616_, _03574_);
    and _10162_(_03618_, _03617_, _03612_);
    or _10163_(_03619_, _03531_, modulus[1]);
    or _10164_(_03620_, _03537_, modulus[0]);
    or _10165_(_03622_, _03620_, _03532_);
    and _10166_(_03623_, _03622_, _03619_);
    and _10167_(_03624_, _03550_, _03546_);
    or _10168_(_03625_, _03624_, _03539_);
    and _10169_(_03626_, _03625_, _03623_);
    or _10170_(_03627_, _03626_, _03575_);
    and _10171_(_03628_, _03627_, _03618_);
    nor _10172_(_03629_, _03591_, _03586_);
    and _10173_(_03630_, _03602_, _03597_);
    or _10174_(_03631_, _03630_, _03592_);
    and _10175_(_03633_, _03631_, _03629_);
    nand _10176_(_03634_, _03604_, _03376_);
    nand _10177_(_03635_, _03634_, _03633_);
    nand _10178_(_03636_, _03635_, _03576_);
    nand _10179_(_03637_, _03636_, _03628_);
    and _10180_(_03638_, _03637_, _00587_);
    nand _10181_(_03639_, _03638_, _06071_);
    nand _10182_(_03640_, _03639_, _03607_);
    or _10183_(_03641_, _03640_, _03524_);
    and _10184_(_03642_, _03634_, _03633_);
    or _10185_(_03644_, _03642_, _03552_);
    and _10186_(_03645_, _03644_, _03626_);
    or _10187_(_03646_, _03645_, _03567_);
    and _10188_(_03647_, _03646_, _03616_);
    or _10189_(_03648_, _03647_, _03573_);
    and _10190_(_03649_, _03648_, _03609_);
    xor _10191_(_03650_, _03649_, _03568_);
    nand _10192_(_03651_, _03650_, _03640_);
    and _10193_(_03652_, _03651_, _03641_);
    or _10194_(_03653_, _03640_, _03531_);
    or _10195_(_03655_, _03642_, _03551_);
    and _10196_(_03656_, _03655_, _03624_);
    or _10197_(_03657_, _03656_, _03538_);
    and _10198_(_03658_, _03657_, _03620_);
    xor _10199_(_03659_, _03658_, _03532_);
    nand _10200_(_03660_, _03659_, _03640_);
    and _10201_(_03661_, _03660_, _03653_);
    xor _10202_(_03662_, _03661_, _00183_);
    or _10203_(_03663_, _03640_, _03537_);
    xor _10204_(_03664_, _03656_, _03538_);
    nand _10205_(_03666_, _03664_, _03640_);
    and _10206_(_03667_, _03666_, _03663_);
    xor _10207_(_03668_, _03667_, _06035_);
    or _10208_(_03669_, _03668_, _03662_);
    or _10209_(_03670_, _03640_, _03546_);
    and _10210_(_03671_, _03639_, _03607_);
    and _10211_(_03672_, _03642_, _03550_);
    xor _10212_(_03673_, _03672_, _03546_);
    or _10213_(_03674_, _03673_, _03671_);
    and _10214_(_03675_, _03674_, _03670_);
    xor _10215_(_03677_, _03675_, _05927_);
    or _10216_(_03678_, _03640_, _03550_);
    xor _10217_(_03679_, _03642_, _03550_);
    or _10218_(_03680_, _03679_, _03671_);
    and _10219_(_03681_, _03680_, _03678_);
    not _10220_(_03682_, _03681_);
    or _10221_(_03683_, _03682_, _03677_);
    or _10222_(_03684_, _03683_, _03669_);
    or _10223_(_03685_, _03640_, _03559_);
    or _10224_(_03686_, _03645_, _03565_);
    and _10225_(_03688_, _03686_, _03614_);
    xor _10226_(_03689_, _03688_, _03560_);
    nand _10227_(_03690_, _03689_, _03640_);
    and _10228_(_03691_, _03690_, _03685_);
    xor _10229_(_03692_, _03691_, _00429_);
    or _10230_(_03693_, _03640_, _03564_);
    xor _10231_(_03694_, _03645_, _03565_);
    nand _10232_(_03695_, _03694_, _03640_);
    and _10233_(_03696_, _03695_, _03693_);
    xor _10234_(_03697_, _03696_, _00309_);
    or _10235_(_03699_, _03697_, _03692_);
    xor _10236_(_03700_, _03652_, _00673_);
    or _10237_(_03701_, _03640_, _03572_);
    xor _10238_(_03702_, _03647_, _03573_);
    nand _10239_(_03703_, _03702_, _03640_);
    and _10240_(_03704_, _03703_, _03701_);
    xor _10241_(_03705_, _03704_, _00550_);
    or _10242_(_03706_, _03705_, _03700_);
    or _10243_(_03707_, _03706_, _03699_);
    nor _10244_(_03708_, _03707_, _03684_);
    not _10245_(_03710_, _03586_);
    or _10246_(_03711_, _03640_, _03710_);
    not _10247_(_03712_, _03591_);
    or _10248_(_03713_, _03603_, _03127_);
    and _10249_(_03714_, _03713_, _03630_);
    and _10250_(_03715_, _03714_, _03712_);
    xor _10251_(_03716_, _03715_, _03710_);
    or _10252_(_03717_, _03716_, _03671_);
    and _10253_(_03718_, _03717_, _03711_);
    or _10254_(_03719_, _03640_, _03712_);
    xor _10255_(_03721_, _03714_, _03712_);
    or _10256_(_03722_, _03721_, _03671_);
    and _10257_(_03723_, _03722_, _03719_);
    nand _10258_(_03724_, _03723_, _03718_);
    or _10259_(_03725_, _03640_, _03597_);
    and _10260_(_03726_, _03602_, _03127_);
    xor _10261_(_03727_, _03726_, _03597_);
    or _10262_(_03728_, _03727_, _03671_);
    and _10263_(_03729_, _03728_, _03725_);
    or _10264_(_03730_, _03640_, _03602_);
    xor _10265_(_03732_, _03602_, _03127_);
    or _10266_(_03733_, _03732_, _03671_);
    and _10267_(_03734_, _03733_, _03730_);
    nand _10268_(_03735_, _03734_, _03729_);
    nor _10269_(_03736_, _03735_, _03724_);
    and _10270_(_03737_, _03736_, _02989_);
    and _10271_(_03738_, _03737_, _03708_);
    nand _10272_(_03739_, _03738_, _00709_);
    or _10273_(_03740_, _03652_, modulus[6]);
    or _10274_(_03741_, _03704_, modulus[5]);
    or _10275_(_03743_, _03741_, _03700_);
    and _10276_(_03744_, _03743_, _03740_);
    or _10277_(_03745_, _03691_, modulus[4]);
    or _10278_(_03746_, _03696_, modulus[3]);
    or _10279_(_03747_, _03746_, _03692_);
    and _10280_(_03748_, _03747_, _03745_);
    or _10281_(_03749_, _03748_, _03706_);
    and _10282_(_03750_, _03749_, _03744_);
    or _10283_(_03751_, _03661_, modulus[2]);
    or _10284_(_03752_, _03667_, modulus[1]);
    or _10285_(_03754_, _03752_, _03662_);
    and _10286_(_03755_, _03754_, _03751_);
    or _10287_(_03756_, _03675_, modulus[0]);
    or _10288_(_03757_, _03681_, _03677_);
    and _10289_(_03758_, _03757_, _03756_);
    or _10290_(_03759_, _03758_, _03669_);
    and _10291_(_03760_, _03759_, _03755_);
    or _10292_(_03761_, _03760_, _03707_);
    and _10293_(_03762_, _03761_, _03750_);
    and _10294_(_03763_, _03723_, _03718_);
    and _10295_(_03765_, _03734_, _03729_);
    or _10296_(_03766_, _03765_, _03724_);
    and _10297_(_03767_, _03766_, _03763_);
    nand _10298_(_03768_, _03736_, _03376_);
    and _10299_(_03769_, _03768_, _03767_);
    not _10300_(_03770_, _03769_);
    nand _10301_(_03771_, _03770_, _03708_);
    nand _10302_(_03772_, _03771_, _03762_);
    and _10303_(_03773_, _03772_, _00708_);
    nand _10304_(_03774_, _03773_, _05956_);
    nand _10305_(_03776_, _03774_, _03739_);
    or _10306_(_03777_, _03776_, _03652_);
    or _10307_(_03778_, _03769_, _03684_);
    and _10308_(_03779_, _03778_, _03760_);
    or _10309_(_03780_, _03779_, _03699_);
    and _10310_(_03781_, _03780_, _03748_);
    or _10311_(_03782_, _03781_, _03705_);
    and _10312_(_03783_, _03782_, _03741_);
    xor _10313_(_03784_, _03783_, _03700_);
    nand _10314_(_03785_, _03784_, _03776_);
    and _10315_(_03787_, _03785_, _03777_);
    or _10316_(_03788_, _03776_, _03661_);
    or _10317_(_03789_, _03769_, _03683_);
    and _10318_(_03790_, _03789_, _03758_);
    or _10319_(_03791_, _03790_, _03668_);
    and _10320_(_03792_, _03791_, _03752_);
    xor _10321_(_03793_, _03792_, _03662_);
    nand _10322_(_03794_, _03793_, _03776_);
    and _10323_(_03795_, _03794_, _03788_);
    xor _10324_(_03796_, _03795_, _00309_);
    or _10325_(_03798_, _03776_, _03667_);
    and _10326_(_03799_, _03774_, _03739_);
    xnor _10327_(_03800_, _03790_, _03668_);
    or _10328_(_03801_, _03800_, _03799_);
    and _10329_(_03802_, _03801_, _03798_);
    xor _10330_(_03803_, _03802_, _00183_);
    or _10331_(_03804_, _03803_, _03796_);
    or _10332_(_03805_, _03776_, _03675_);
    and _10333_(_03806_, _03769_, _03681_);
    xnor _10334_(_03807_, _03806_, _03677_);
    or _10335_(_03809_, _03807_, _03799_);
    and _10336_(_03810_, _03809_, _03805_);
    xor _10337_(_03811_, _03810_, _06035_);
    or _10338_(_03812_, _03776_, _03681_);
    xor _10339_(_03813_, _03769_, _03681_);
    or _10340_(_03814_, _03813_, _03799_);
    and _10341_(_03815_, _03814_, _03812_);
    xor _10342_(_03816_, _03815_, _05927_);
    or _10343_(_03817_, _03816_, _03811_);
    or _10344_(_03818_, _03817_, _03804_);
    or _10345_(_03820_, _03776_, _03691_);
    or _10346_(_03821_, _03779_, _03697_);
    and _10347_(_03822_, _03821_, _03746_);
    xor _10348_(_03823_, _03822_, _03692_);
    nand _10349_(_03824_, _03823_, _03776_);
    and _10350_(_03825_, _03824_, _03820_);
    xor _10351_(_03826_, _03825_, _00550_);
    or _10352_(_03827_, _03776_, _03696_);
    xnor _10353_(_03828_, _03779_, _03697_);
    or _10354_(_03829_, _03828_, _03799_);
    and _10355_(_03831_, _03829_, _03827_);
    xor _10356_(_03832_, _03831_, _00429_);
    or _10357_(_03833_, _03832_, _03826_);
    xor _10358_(_03834_, _03787_, _00797_);
    or _10359_(_03835_, _03776_, _03704_);
    xor _10360_(_03836_, _03781_, _03705_);
    nand _10361_(_03837_, _03836_, _03776_);
    and _10362_(_03838_, _03837_, _03835_);
    xor _10363_(_03839_, _03838_, _00673_);
    or _10364_(_03840_, _03839_, _03834_);
    or _10365_(_03842_, _03840_, _03833_);
    nor _10366_(_03843_, _03842_, _03818_);
    or _10367_(_03844_, _03776_, _03718_);
    or _10368_(_03845_, _03735_, _03127_);
    and _10369_(_03846_, _03845_, _03765_);
    and _10370_(_03847_, _03846_, _03723_);
    xor _10371_(_03848_, _03847_, _03718_);
    or _10372_(_03849_, _03848_, _03799_);
    nand _10373_(_03850_, _03849_, _03844_);
    or _10374_(_03851_, _03776_, _03723_);
    xor _10375_(_03853_, _03846_, _03723_);
    or _10376_(_03854_, _03853_, _03799_);
    nand _10377_(_03855_, _03854_, _03851_);
    or _10378_(_03856_, _03855_, _03850_);
    or _10379_(_03857_, _03776_, _03729_);
    and _10380_(_03858_, _03734_, _03127_);
    xor _10381_(_03859_, _03858_, _03729_);
    or _10382_(_03860_, _03859_, _03799_);
    and _10383_(_03861_, _03860_, _03857_);
    or _10384_(_03862_, _03776_, _03734_);
    xor _10385_(_03864_, _03734_, _03127_);
    or _10386_(_03865_, _03864_, _03799_);
    and _10387_(_03866_, _03865_, _03862_);
    nand _10388_(_03867_, _03866_, _03861_);
    nor _10389_(_03868_, _03867_, _03856_);
    and _10390_(_03869_, _03868_, _02989_);
    and _10391_(_03870_, _03869_, _03843_);
    nand _10392_(_03871_, _03870_, _00754_);
    or _10393_(_03872_, _03787_, modulus[7]);
    or _10394_(_03873_, _03838_, modulus[6]);
    or _10395_(_03875_, _03873_, _03834_);
    and _10396_(_03876_, _03875_, _03872_);
    or _10397_(_03877_, _03825_, modulus[5]);
    or _10398_(_03878_, _03831_, modulus[4]);
    or _10399_(_03879_, _03878_, _03826_);
    and _10400_(_03880_, _03879_, _03877_);
    or _10401_(_03881_, _03880_, _03840_);
    and _10402_(_03882_, _03881_, _03876_);
    or _10403_(_03883_, _03795_, modulus[3]);
    or _10404_(_03884_, _03802_, modulus[2]);
    or _10405_(_03886_, _03884_, _03796_);
    and _10406_(_03887_, _03886_, _03883_);
    or _10407_(_03888_, _03810_, modulus[1]);
    or _10408_(_03889_, _03815_, modulus[0]);
    or _10409_(_03890_, _03889_, _03811_);
    and _10410_(_03891_, _03890_, _03888_);
    or _10411_(_03892_, _03891_, _03804_);
    and _10412_(_03893_, _03892_, _03887_);
    or _10413_(_03894_, _03893_, _03842_);
    and _10414_(_03895_, _03894_, _03882_);
    nor _10415_(_03897_, _03855_, _03850_);
    and _10416_(_03898_, _03866_, _03861_);
    or _10417_(_03899_, _03898_, _03856_);
    and _10418_(_03900_, _03899_, _03897_);
    nand _10419_(_03901_, _03868_, _03376_);
    and _10420_(_03902_, _03901_, _03900_);
    not _10421_(_03903_, _03902_);
    nand _10422_(_03904_, _03903_, _03843_);
    nand _10423_(_03905_, _03904_, _03895_);
    nand _10424_(_03906_, _03905_, _00754_);
    nand _10425_(_03908_, _03906_, _03871_);
    or _10426_(_03909_, _03908_, _03787_);
    or _10427_(_03910_, _03902_, _03818_);
    and _10428_(_03911_, _03910_, _03893_);
    or _10429_(_03912_, _03911_, _03833_);
    and _10430_(_03913_, _03912_, _03880_);
    or _10431_(_03914_, _03913_, _03839_);
    and _10432_(_03915_, _03914_, _03873_);
    xor _10433_(_03916_, _03915_, _03834_);
    nand _10434_(_03917_, _03916_, _03908_);
    and _10435_(_03919_, _03917_, _03909_);
    or _10436_(_03920_, _03908_, _03795_);
    or _10437_(_03921_, _03902_, _03817_);
    and _10438_(_03922_, _03921_, _03891_);
    or _10439_(_03923_, _03922_, _03803_);
    and _10440_(_03924_, _03923_, _03884_);
    xor _10441_(_03925_, _03924_, _03796_);
    nand _10442_(_03926_, _03925_, _03908_);
    and _10443_(_03927_, _03926_, _03920_);
    xor _10444_(_03928_, _03927_, _00429_);
    or _10445_(_03930_, _03908_, _03802_);
    xor _10446_(_03931_, _03922_, _03803_);
    nand _10447_(_03932_, _03931_, _03908_);
    and _10448_(_03933_, _03932_, _03930_);
    xor _10449_(_03934_, _03933_, _00309_);
    or _10450_(_03935_, _03934_, _03928_);
    or _10451_(_03936_, _03908_, _03810_);
    or _10452_(_03937_, _03902_, _03816_);
    and _10453_(_03938_, _03937_, _03889_);
    xor _10454_(_03939_, _03938_, _03811_);
    nand _10455_(_03941_, _03939_, _03908_);
    and _10456_(_03942_, _03941_, _03936_);
    xor _10457_(_03943_, _03942_, _00183_);
    or _10458_(_03944_, _03908_, _03815_);
    and _10459_(_03945_, _03906_, _03871_);
    xnor _10460_(_03946_, _03902_, _03816_);
    or _10461_(_03947_, _03946_, _03945_);
    and _10462_(_03948_, _03947_, _03944_);
    xor _10463_(_03949_, _03948_, _06035_);
    or _10464_(_03950_, _03949_, _03943_);
    or _10465_(_03952_, _03950_, _03935_);
    or _10466_(_03953_, _03908_, _03825_);
    or _10467_(_03954_, _03911_, _03832_);
    and _10468_(_03955_, _03954_, _03878_);
    xor _10469_(_03956_, _03955_, _03826_);
    nand _10470_(_03957_, _03956_, _03908_);
    and _10471_(_03958_, _03957_, _03953_);
    xor _10472_(_03959_, _03958_, _00673_);
    or _10473_(_03960_, _03908_, _03831_);
    xor _10474_(_03961_, _03911_, _03832_);
    nand _10475_(_03963_, _03961_, _03908_);
    and _10476_(_03964_, _03963_, _03960_);
    xor _10477_(_03965_, _03964_, _00550_);
    or _10478_(_03966_, _03965_, _03959_);
    xor _10479_(_03967_, _03919_, _00919_);
    or _10480_(_03968_, _03908_, _03838_);
    xor _10481_(_03969_, _03913_, _03839_);
    nand _10482_(_03970_, _03969_, _03908_);
    and _10483_(_03971_, _03970_, _03968_);
    xor _10484_(_03972_, _03971_, _00797_);
    or _10485_(_03974_, _03972_, _03967_);
    or _10486_(_03975_, _03974_, _03966_);
    nor _10487_(_03976_, _03975_, _03952_);
    not _10488_(_03977_, _03850_);
    or _10489_(_03978_, _03908_, _03977_);
    not _10490_(_03979_, _03855_);
    or _10491_(_03980_, _03867_, _03127_);
    and _10492_(_03981_, _03980_, _03898_);
    and _10493_(_03982_, _03981_, _03979_);
    xor _10494_(_03983_, _03982_, _03977_);
    or _10495_(_03985_, _03983_, _03945_);
    and _10496_(_03986_, _03985_, _03978_);
    xor _10497_(_03987_, _03986_, _05927_);
    or _10498_(_03988_, _03908_, _03979_);
    xor _10499_(_03989_, _03981_, _03979_);
    or _10500_(_03990_, _03989_, _03945_);
    and _10501_(_03991_, _03990_, _03988_);
    not _10502_(_03992_, _03991_);
    or _10503_(_03993_, _03992_, _03987_);
    or _10504_(_03994_, _03908_, _03861_);
    and _10505_(_03996_, _03866_, _03127_);
    xor _10506_(_03997_, _03996_, _03861_);
    or _10507_(_03998_, _03997_, _03945_);
    and _10508_(_03999_, _03998_, _03994_);
    or _10509_(_04000_, _03908_, _03866_);
    xor _10510_(_04001_, _03866_, _03127_);
    or _10511_(_04002_, _04001_, _03945_);
    and _10512_(_04003_, _04002_, _04000_);
    nand _10513_(_04004_, _04003_, _03999_);
    nor _10514_(_04005_, _04004_, _03993_);
    and _10515_(_04007_, _04005_, _02989_);
    and _10516_(_04008_, _04007_, _03976_);
    nand _10517_(_04009_, _04008_, _05959_);
    or _10518_(_04010_, _03919_, modulus[8]);
    or _10519_(_04011_, _03971_, modulus[7]);
    or _10520_(_04012_, _04011_, _03967_);
    and _10521_(_04013_, _04012_, _04010_);
    or _10522_(_04014_, _03958_, modulus[6]);
    or _10523_(_04015_, _03964_, modulus[5]);
    or _10524_(_04016_, _04015_, _03959_);
    and _10525_(_04018_, _04016_, _04014_);
    or _10526_(_04019_, _04018_, _03974_);
    and _10527_(_04020_, _04019_, _04013_);
    or _10528_(_04021_, _03927_, modulus[4]);
    or _10529_(_04022_, _03933_, modulus[3]);
    or _10530_(_04023_, _04022_, _03928_);
    and _10531_(_04024_, _04023_, _04021_);
    or _10532_(_04025_, _03942_, modulus[2]);
    or _10533_(_04026_, _03948_, modulus[1]);
    or _10534_(_04027_, _04026_, _03943_);
    and _10535_(_04029_, _04027_, _04025_);
    or _10536_(_04030_, _04029_, _03935_);
    and _10537_(_04031_, _04030_, _04024_);
    or _10538_(_04032_, _04031_, _03975_);
    and _10539_(_04033_, _04032_, _04020_);
    or _10540_(_04034_, _03986_, modulus[0]);
    or _10541_(_04035_, _03991_, _03987_);
    and _10542_(_04036_, _04035_, _04034_);
    and _10543_(_04037_, _04003_, _03999_);
    or _10544_(_04038_, _04037_, _03993_);
    and _10545_(_04040_, _04038_, _04036_);
    nand _10546_(_04041_, _04005_, _03376_);
    nand _10547_(_04042_, _04041_, _04040_);
    nand _10548_(_04043_, _04042_, _03976_);
    nand _10549_(_04044_, _04043_, _04033_);
    and _10550_(_04045_, _04044_, _05955_);
    and _10551_(_04046_, _04045_, _05957_);
    nand _10552_(_04047_, _04046_, _05956_);
    nand _10553_(_04048_, _04047_, _04009_);
    or _10554_(_04049_, _04048_, _03919_);
    not _10555_(_04051_, _04042_);
    or _10556_(_04052_, _04051_, _03952_);
    and _10557_(_04053_, _04052_, _04031_);
    or _10558_(_04054_, _04053_, _03966_);
    and _10559_(_04055_, _04054_, _04018_);
    or _10560_(_04056_, _04055_, _03972_);
    and _10561_(_04057_, _04056_, _04011_);
    xor _10562_(_04058_, _04057_, _03967_);
    nand _10563_(_04059_, _04058_, _04048_);
    and _10564_(_04060_, _04059_, _04049_);
    or _10565_(_04062_, _04048_, _03927_);
    or _10566_(_04063_, _04051_, _03950_);
    and _10567_(_04064_, _04063_, _04029_);
    or _10568_(_04065_, _04064_, _03934_);
    and _10569_(_04066_, _04065_, _04022_);
    xor _10570_(_04067_, _04066_, _03928_);
    nand _10571_(_04068_, _04067_, _04048_);
    and _10572_(_04069_, _04068_, _04062_);
    xor _10573_(_04070_, _04069_, _00550_);
    or _10574_(_04071_, _04048_, _03933_);
    and _10575_(_04073_, _04047_, _04009_);
    xnor _10576_(_04074_, _04064_, _03934_);
    or _10577_(_04075_, _04074_, _04073_);
    and _10578_(_04076_, _04075_, _04071_);
    xor _10579_(_04077_, _04076_, _00429_);
    or _10580_(_04078_, _04077_, _04070_);
    or _10581_(_04079_, _04048_, _03942_);
    or _10582_(_04080_, _04051_, _03949_);
    and _10583_(_04081_, _04080_, _04026_);
    xnor _10584_(_04082_, _04081_, _03943_);
    or _10585_(_04084_, _04082_, _04073_);
    and _10586_(_04085_, _04084_, _04079_);
    xor _10587_(_04086_, _04085_, _00309_);
    or _10588_(_04087_, _04048_, _03948_);
    xor _10589_(_04088_, _04042_, _03949_);
    or _10590_(_04089_, _04088_, _04073_);
    and _10591_(_04090_, _04089_, _04087_);
    xor _10592_(_04091_, _04090_, _00183_);
    or _10593_(_04092_, _04091_, _04086_);
    or _10594_(_04093_, _04092_, _04078_);
    or _10595_(_04095_, _04048_, _03958_);
    or _10596_(_04096_, _04053_, _03965_);
    and _10597_(_04097_, _04096_, _04015_);
    xor _10598_(_04098_, _04097_, _03959_);
    nand _10599_(_04099_, _04098_, _04048_);
    and _10600_(_04100_, _04099_, _04095_);
    xor _10601_(_04101_, _04100_, _00797_);
    or _10602_(_04102_, _04048_, _03964_);
    xnor _10603_(_04103_, _04053_, _03965_);
    or _10604_(_04104_, _04103_, _04073_);
    and _10605_(_04106_, _04104_, _04102_);
    xor _10606_(_04107_, _04106_, _00673_);
    or _10607_(_04108_, _04107_, _04101_);
    xor _10608_(_04109_, _04060_, _01048_);
    or _10609_(_04110_, _04048_, _03971_);
    xor _10610_(_04111_, _04055_, _03972_);
    nand _10611_(_04112_, _04111_, _04048_);
    and _10612_(_04113_, _04112_, _04110_);
    xor _10613_(_04114_, _04113_, _00919_);
    or _10614_(_04115_, _04114_, _04109_);
    or _10615_(_04117_, _04115_, _04108_);
    nor _10616_(_04118_, _04117_, _04093_);
    or _10617_(_04119_, _04048_, _03986_);
    or _10618_(_04120_, _04004_, _03127_);
    and _10619_(_04121_, _04120_, _04037_);
    and _10620_(_04122_, _04121_, _03991_);
    xnor _10621_(_04123_, _04122_, _03987_);
    or _10622_(_04124_, _04123_, _04073_);
    and _10623_(_04125_, _04124_, _04119_);
    xor _10624_(_04126_, _04125_, _06035_);
    or _10625_(_04128_, _04048_, _03991_);
    xor _10626_(_04129_, _04121_, _03991_);
    or _10627_(_04130_, _04129_, _04073_);
    and _10628_(_04131_, _04130_, _04128_);
    xor _10629_(_04132_, _04131_, _05927_);
    or _10630_(_04133_, _04132_, _04126_);
    or _10631_(_04134_, _04048_, _03999_);
    and _10632_(_04135_, _04003_, _03127_);
    xor _10633_(_04136_, _04135_, _03999_);
    or _10634_(_04137_, _04136_, _04073_);
    and _10635_(_04139_, _04137_, _04134_);
    or _10636_(_04140_, _04048_, _04003_);
    xor _10637_(_04141_, _04003_, _03127_);
    or _10638_(_04142_, _04141_, _04073_);
    and _10639_(_04143_, _04142_, _04140_);
    nand _10640_(_04144_, _04143_, _04139_);
    nor _10641_(_04145_, _04144_, _04133_);
    and _10642_(_04146_, _04145_, _02989_);
    and _10643_(_04147_, _04146_, _04118_);
    nand _10644_(_04148_, _04147_, _06075_);
    or _10645_(_04150_, _04060_, modulus[9]);
    or _10646_(_04151_, _04113_, modulus[8]);
    or _10647_(_04152_, _04151_, _04109_);
    and _10648_(_04153_, _04152_, _04150_);
    or _10649_(_04154_, _04100_, modulus[7]);
    or _10650_(_04155_, _04106_, modulus[6]);
    or _10651_(_04156_, _04155_, _04101_);
    and _10652_(_04157_, _04156_, _04154_);
    or _10653_(_04158_, _04157_, _04115_);
    and _10654_(_04159_, _04158_, _04153_);
    or _10655_(_04161_, _04069_, modulus[5]);
    or _10656_(_04162_, _04076_, modulus[4]);
    or _10657_(_04163_, _04162_, _04070_);
    and _10658_(_04164_, _04163_, _04161_);
    or _10659_(_04165_, _04085_, modulus[3]);
    or _10660_(_04166_, _04090_, modulus[2]);
    or _10661_(_04167_, _04166_, _04086_);
    and _10662_(_04168_, _04167_, _04165_);
    or _10663_(_04169_, _04168_, _04078_);
    and _10664_(_04170_, _04169_, _04164_);
    or _10665_(_04172_, _04170_, _04117_);
    and _10666_(_04173_, _04172_, _04159_);
    or _10667_(_04174_, _04125_, modulus[1]);
    or _10668_(_04175_, _04131_, modulus[0]);
    or _10669_(_04176_, _04175_, _04126_);
    and _10670_(_04177_, _04176_, _04174_);
    and _10671_(_04178_, _04143_, _04139_);
    or _10672_(_04179_, _04178_, _04133_);
    and _10673_(_04180_, _04179_, _04177_);
    nand _10674_(_04181_, _04145_, _03376_);
    nand _10675_(_04183_, _04181_, _04180_);
    nand _10676_(_04184_, _04183_, _04118_);
    nand _10677_(_04185_, _04184_, _04173_);
    and _10678_(_04186_, _04185_, _06074_);
    nand _10679_(_04187_, _04186_, _06071_);
    nand _10680_(_04188_, _04187_, _04148_);
    or _10681_(_04189_, _04188_, _04060_);
    and _10682_(_04190_, _04181_, _04180_);
    or _10683_(_04191_, _04190_, _04093_);
    and _10684_(_04192_, _04191_, _04170_);
    or _10685_(_04194_, _04192_, _04108_);
    and _10686_(_04195_, _04194_, _04157_);
    or _10687_(_04196_, _04195_, _04114_);
    and _10688_(_04197_, _04196_, _04151_);
    xor _10689_(_04198_, _04197_, _04109_);
    nand _10690_(_04199_, _04198_, _04188_);
    and _10691_(_04200_, _04199_, _04189_);
    or _10692_(_04201_, _04188_, _04069_);
    or _10693_(_04202_, _04190_, _04092_);
    and _10694_(_04203_, _04202_, _04168_);
    or _10695_(_04205_, _04203_, _04077_);
    and _10696_(_04206_, _04205_, _04162_);
    xor _10697_(_04207_, _04206_, _04070_);
    nand _10698_(_04208_, _04207_, _04188_);
    and _10699_(_04209_, _04208_, _04201_);
    xor _10700_(_04210_, _04209_, _00673_);
    or _10701_(_04211_, _04188_, _04076_);
    xor _10702_(_04212_, _04203_, _04077_);
    nand _10703_(_04213_, _04212_, _04188_);
    and _10704_(_04214_, _04213_, _04211_);
    xor _10705_(_04216_, _04214_, _00550_);
    or _10706_(_04217_, _04216_, _04210_);
    or _10707_(_04218_, _04188_, _04085_);
    or _10708_(_04219_, _04190_, _04091_);
    and _10709_(_04220_, _04219_, _04166_);
    xor _10710_(_04221_, _04220_, _04086_);
    nand _10711_(_04222_, _04221_, _04188_);
    and _10712_(_04223_, _04222_, _04218_);
    xor _10713_(_04224_, _04223_, _00429_);
    or _10714_(_04225_, _04188_, _04090_);
    and _10715_(_04227_, _04187_, _04148_);
    xor _10716_(_04228_, _04183_, _04091_);
    or _10717_(_04229_, _04228_, _04227_);
    and _10718_(_04230_, _04229_, _04225_);
    xor _10719_(_04231_, _04230_, _00309_);
    or _10720_(_04232_, _04231_, _04224_);
    or _10721_(_04233_, _04232_, _04217_);
    or _10722_(_04234_, _04188_, _04100_);
    or _10723_(_04235_, _04192_, _04107_);
    and _10724_(_04236_, _04235_, _04155_);
    xor _10725_(_04238_, _04236_, _04101_);
    nand _10726_(_04239_, _04238_, _04188_);
    and _10727_(_04240_, _04239_, _04234_);
    xor _10728_(_04241_, _04240_, _00919_);
    or _10729_(_04242_, _04188_, _04106_);
    xor _10730_(_04243_, _04192_, _04107_);
    nand _10731_(_04244_, _04243_, _04188_);
    and _10732_(_04245_, _04244_, _04242_);
    xor _10733_(_04246_, _04245_, _00797_);
    or _10734_(_04247_, _04246_, _04241_);
    xor _10735_(_04249_, _04200_, _01181_);
    or _10736_(_04250_, _04188_, _04113_);
    xor _10737_(_04251_, _04195_, _04114_);
    nand _10738_(_04252_, _04251_, _04188_);
    and _10739_(_04253_, _04252_, _04250_);
    xor _10740_(_04254_, _04253_, _01048_);
    or _10741_(_04255_, _04254_, _04249_);
    or _10742_(_04256_, _04255_, _04247_);
    nor _10743_(_04257_, _04256_, _04233_);
    or _10744_(_04258_, _04188_, _04125_);
    or _10745_(_04260_, _04144_, _03127_);
    and _10746_(_04261_, _04260_, _04178_);
    or _10747_(_04262_, _04261_, _04132_);
    and _10748_(_04263_, _04262_, _04175_);
    xnor _10749_(_04264_, _04263_, _04126_);
    or _10750_(_04265_, _04264_, _04227_);
    and _10751_(_04266_, _04265_, _04258_);
    xor _10752_(_04267_, _04266_, _00183_);
    or _10753_(_04268_, _04188_, _04131_);
    xnor _10754_(_04269_, _04261_, _04132_);
    or _10755_(_04271_, _04269_, _04227_);
    and _10756_(_04272_, _04271_, _04268_);
    xor _10757_(_04273_, _04272_, _06035_);
    or _10758_(_04274_, _04273_, _04267_);
    or _10759_(_04275_, _04188_, _04139_);
    and _10760_(_04276_, _04143_, _03127_);
    xor _10761_(_04277_, _04276_, _04139_);
    or _10762_(_04278_, _04277_, _04227_);
    and _10763_(_04279_, _04278_, _04275_);
    xor _10764_(_04280_, _04279_, _05927_);
    or _10765_(_04282_, _04188_, _04143_);
    xor _10766_(_04283_, _04143_, _03127_);
    or _10767_(_04284_, _04283_, _04227_);
    and _10768_(_04285_, _04284_, _04282_);
    not _10769_(_04286_, _04285_);
    or _10770_(_04287_, _04286_, _04280_);
    nor _10771_(_04288_, _04287_, _04274_);
    and _10772_(_04289_, _04288_, _02989_);
    and _10773_(_04290_, _04289_, _04257_);
    nand _10774_(_04291_, _04290_, _00230_);
    or _10775_(_04293_, _04200_, modulus[10]);
    or _10776_(_04294_, _04253_, modulus[9]);
    or _10777_(_04295_, _04294_, _04249_);
    and _10778_(_04296_, _04295_, _04293_);
    or _10779_(_04297_, _04240_, modulus[8]);
    or _10780_(_04298_, _04245_, modulus[7]);
    or _10781_(_04299_, _04298_, _04241_);
    and _10782_(_04300_, _04299_, _04297_);
    or _10783_(_04301_, _04300_, _04255_);
    and _10784_(_04302_, _04301_, _04296_);
    or _10785_(_04304_, _04209_, modulus[6]);
    or _10786_(_04305_, _04214_, modulus[5]);
    or _10787_(_04306_, _04305_, _04210_);
    and _10788_(_04307_, _04306_, _04304_);
    or _10789_(_04308_, _04223_, modulus[4]);
    or _10790_(_04309_, _04230_, modulus[3]);
    or _10791_(_04310_, _04309_, _04224_);
    and _10792_(_04311_, _04310_, _04308_);
    or _10793_(_04312_, _04311_, _04217_);
    and _10794_(_04313_, _04312_, _04307_);
    or _10795_(_04315_, _04313_, _04256_);
    and _10796_(_04316_, _04315_, _04302_);
    or _10797_(_04317_, _04266_, modulus[2]);
    or _10798_(_04318_, _04272_, modulus[1]);
    or _10799_(_04319_, _04318_, _04267_);
    and _10800_(_04320_, _04319_, _04317_);
    or _10801_(_04321_, _04279_, modulus[0]);
    or _10802_(_04322_, _04285_, _04280_);
    and _10803_(_04323_, _04322_, _04321_);
    or _10804_(_04324_, _04323_, _04274_);
    and _10805_(_04326_, _04324_, _04320_);
    nand _10806_(_04327_, _04288_, _03376_);
    nand _10807_(_04328_, _04327_, _04326_);
    nand _10808_(_04329_, _04328_, _04257_);
    nand _10809_(_04330_, _04329_, _04316_);
    and _10810_(_04331_, _04330_, _00229_);
    nand _10811_(_04332_, _04331_, _05956_);
    nand _10812_(_04333_, _04332_, _04291_);
    or _10813_(_04334_, _04333_, _04200_);
    and _10814_(_04335_, _04327_, _04326_);
    or _10815_(_04337_, _04335_, _04233_);
    and _10816_(_04338_, _04337_, _04313_);
    or _10817_(_04339_, _04338_, _04247_);
    and _10818_(_04340_, _04339_, _04300_);
    or _10819_(_04341_, _04340_, _04254_);
    and _10820_(_04342_, _04341_, _04294_);
    xor _10821_(_04343_, _04342_, _04249_);
    nand _10822_(_04344_, _04343_, _04333_);
    and _10823_(_04345_, _04344_, _04334_);
    or _10824_(_04346_, _04333_, _04209_);
    or _10825_(_04348_, _04335_, _04232_);
    and _10826_(_04349_, _04348_, _04311_);
    or _10827_(_04350_, _04349_, _04216_);
    and _10828_(_04351_, _04350_, _04305_);
    xor _10829_(_04352_, _04351_, _04210_);
    nand _10830_(_04353_, _04352_, _04333_);
    and _10831_(_04354_, _04353_, _04346_);
    xor _10832_(_04355_, _04354_, _00797_);
    or _10833_(_04356_, _04333_, _04214_);
    xor _10834_(_04357_, _04349_, _04216_);
    nand _10835_(_04359_, _04357_, _04333_);
    and _10836_(_04360_, _04359_, _04356_);
    xor _10837_(_04361_, _04360_, _00673_);
    or _10838_(_04362_, _04361_, _04355_);
    or _10839_(_04363_, _04333_, _04223_);
    or _10840_(_04364_, _04335_, _04231_);
    and _10841_(_04365_, _04364_, _04309_);
    xor _10842_(_04366_, _04365_, _04224_);
    nand _10843_(_04367_, _04366_, _04333_);
    and _10844_(_04368_, _04367_, _04363_);
    xor _10845_(_04370_, _04368_, _00550_);
    or _10846_(_04371_, _04333_, _04230_);
    and _10847_(_04372_, _04332_, _04291_);
    xor _10848_(_04373_, _04328_, _04231_);
    or _10849_(_04374_, _04373_, _04372_);
    and _10850_(_04375_, _04374_, _04371_);
    xor _10851_(_04376_, _04375_, _00429_);
    or _10852_(_04377_, _04376_, _04370_);
    or _10853_(_04378_, _04377_, _04362_);
    or _10854_(_04379_, _04333_, _04240_);
    or _10855_(_04381_, _04338_, _04246_);
    and _10856_(_04382_, _04381_, _04298_);
    xor _10857_(_04383_, _04382_, _04241_);
    nand _10858_(_04384_, _04383_, _04333_);
    and _10859_(_04385_, _04384_, _04379_);
    xor _10860_(_04386_, _04385_, _01048_);
    or _10861_(_04387_, _04333_, _04245_);
    xor _10862_(_04388_, _04338_, _04246_);
    nand _10863_(_04389_, _04388_, _04333_);
    and _10864_(_04390_, _04389_, _04387_);
    xor _10865_(_04392_, _04390_, _00919_);
    or _10866_(_04393_, _04392_, _04386_);
    xor _10867_(_04394_, _04345_, _01328_);
    or _10868_(_04395_, _04333_, _04253_);
    xor _10869_(_04396_, _04340_, _04254_);
    nand _10870_(_04397_, _04396_, _04333_);
    and _10871_(_04398_, _04397_, _04395_);
    xor _10872_(_04399_, _04398_, _01181_);
    or _10873_(_04400_, _04399_, _04394_);
    or _10874_(_04401_, _04400_, _04393_);
    nor _10875_(_04403_, _04401_, _04378_);
    or _10876_(_04404_, _04333_, _04266_);
    or _10877_(_04405_, _04287_, _03127_);
    and _10878_(_04406_, _04405_, _04323_);
    or _10879_(_04407_, _04406_, _04273_);
    and _10880_(_04408_, _04407_, _04318_);
    xnor _10881_(_04409_, _04408_, _04267_);
    or _10882_(_04410_, _04409_, _04372_);
    and _10883_(_04411_, _04410_, _04404_);
    xor _10884_(_04412_, _04411_, _00309_);
    or _10885_(_04414_, _04333_, _04272_);
    xnor _10886_(_04415_, _04406_, _04273_);
    or _10887_(_04416_, _04415_, _04372_);
    and _10888_(_04417_, _04416_, _04414_);
    xor _10889_(_04418_, _04417_, _00183_);
    or _10890_(_04419_, _04418_, _04412_);
    or _10891_(_04420_, _04333_, _04279_);
    and _10892_(_04421_, _04285_, _03127_);
    xnor _10893_(_04422_, _04421_, _04280_);
    or _10894_(_04423_, _04422_, _04372_);
    and _10895_(_04425_, _04423_, _04420_);
    xor _10896_(_04426_, _04425_, _06035_);
    or _10897_(_04427_, _04333_, _04285_);
    xor _10898_(_04428_, _04285_, _03127_);
    or _10899_(_04429_, _04428_, _04372_);
    and _10900_(_04430_, _04429_, _04427_);
    xor _10901_(_04431_, _04430_, _05927_);
    or _10902_(_04432_, _04431_, _04426_);
    nor _10903_(_04433_, _04432_, _04419_);
    and _10904_(_04434_, _04433_, _02989_);
    and _10905_(_04436_, _04434_, _04403_);
    nand _10906_(_04437_, _04436_, _00346_);
    or _10907_(_04438_, _04345_, modulus[11]);
    or _10908_(_04439_, _04398_, modulus[10]);
    or _10909_(_04440_, _04439_, _04394_);
    and _10910_(_04441_, _04440_, _04438_);
    or _10911_(_04442_, _04385_, modulus[9]);
    or _10912_(_04443_, _04390_, modulus[8]);
    or _10913_(_04444_, _04443_, _04386_);
    and _10914_(_04445_, _04444_, _04442_);
    or _10915_(_04447_, _04445_, _04400_);
    and _10916_(_04448_, _04447_, _04441_);
    or _10917_(_04449_, _04354_, modulus[7]);
    or _10918_(_04450_, _04360_, modulus[6]);
    or _10919_(_04451_, _04450_, _04355_);
    and _10920_(_04452_, _04451_, _04449_);
    or _10921_(_04453_, _04368_, modulus[5]);
    or _10922_(_04454_, _04375_, modulus[4]);
    or _10923_(_04455_, _04454_, _04370_);
    and _10924_(_04456_, _04455_, _04453_);
    or _10925_(_04458_, _04456_, _04362_);
    and _10926_(_04459_, _04458_, _04452_);
    or _10927_(_04460_, _04459_, _04401_);
    and _10928_(_04461_, _04460_, _04448_);
    or _10929_(_04462_, _04411_, modulus[3]);
    or _10930_(_04463_, _04417_, modulus[2]);
    or _10931_(_04464_, _04463_, _04412_);
    and _10932_(_04465_, _04464_, _04462_);
    or _10933_(_04466_, _04425_, modulus[1]);
    or _10934_(_04467_, _04430_, modulus[0]);
    or _10935_(_04469_, _04467_, _04426_);
    and _10936_(_04470_, _04469_, _04466_);
    or _10937_(_04471_, _04470_, _04419_);
    and _10938_(_04472_, _04471_, _04465_);
    nand _10939_(_04473_, _04433_, _03376_);
    nand _10940_(_04474_, _04473_, _04472_);
    nand _10941_(_04475_, _04474_, _04403_);
    nand _10942_(_04476_, _04475_, _04461_);
    nand _10943_(_04477_, _04476_, _00346_);
    nand _10944_(_04478_, _04477_, _04437_);
    or _10945_(_04480_, _04478_, _04345_);
    and _10946_(_04481_, _04473_, _04472_);
    or _10947_(_04482_, _04481_, _04378_);
    and _10948_(_04483_, _04482_, _04459_);
    or _10949_(_04484_, _04483_, _04393_);
    and _10950_(_04485_, _04484_, _04445_);
    or _10951_(_04486_, _04485_, _04399_);
    and _10952_(_04487_, _04486_, _04439_);
    xor _10953_(_04488_, _04487_, _04394_);
    nand _10954_(_04489_, _04488_, _04478_);
    and _10955_(_04491_, _04489_, _04480_);
    or _10956_(_04492_, _04478_, _04354_);
    or _10957_(_04493_, _04481_, _04377_);
    and _10958_(_04494_, _04493_, _04456_);
    or _10959_(_04495_, _04494_, _04361_);
    and _10960_(_04496_, _04495_, _04450_);
    xor _10961_(_04497_, _04496_, _04355_);
    nand _10962_(_04498_, _04497_, _04478_);
    and _10963_(_04499_, _04498_, _04492_);
    xor _10964_(_04500_, _04499_, _00919_);
    or _10965_(_04502_, _04478_, _04360_);
    xor _10966_(_04503_, _04494_, _04361_);
    nand _10967_(_04504_, _04503_, _04478_);
    and _10968_(_04505_, _04504_, _04502_);
    xor _10969_(_04506_, _04505_, _00797_);
    or _10970_(_04507_, _04506_, _04500_);
    or _10971_(_04508_, _04478_, _04368_);
    or _10972_(_04509_, _04481_, _04376_);
    and _10973_(_04510_, _04509_, _04454_);
    xor _10974_(_04511_, _04510_, _04370_);
    nand _10975_(_04513_, _04511_, _04478_);
    and _10976_(_04514_, _04513_, _04508_);
    xor _10977_(_04515_, _04514_, _00673_);
    or _10978_(_04516_, _04478_, _04375_);
    xor _10979_(_04517_, _04481_, _04376_);
    nand _10980_(_04518_, _04517_, _04478_);
    and _10981_(_04519_, _04518_, _04516_);
    xor _10982_(_04520_, _04519_, _00550_);
    or _10983_(_04521_, _04520_, _04515_);
    or _10984_(_04522_, _04521_, _04507_);
    or _10985_(_04524_, _04478_, _04385_);
    or _10986_(_04525_, _04483_, _04392_);
    and _10987_(_04526_, _04525_, _04443_);
    xor _10988_(_04527_, _04526_, _04386_);
    nand _10989_(_04528_, _04527_, _04478_);
    and _10990_(_04529_, _04528_, _04524_);
    xor _10991_(_04530_, _04529_, _01181_);
    or _10992_(_04531_, _04478_, _04390_);
    xor _10993_(_04532_, _04483_, _04392_);
    nand _10994_(_04533_, _04532_, _04478_);
    and _10995_(_04535_, _04533_, _04531_);
    xor _10996_(_04536_, _04535_, _01048_);
    or _10997_(_04537_, _04536_, _04530_);
    xor _10998_(_04538_, _04491_, _01474_);
    or _10999_(_04539_, _04478_, _04398_);
    xor _11000_(_04540_, _04485_, _04399_);
    nand _11001_(_04541_, _04540_, _04478_);
    and _11002_(_04542_, _04541_, _04539_);
    xor _11003_(_04543_, _04542_, _01328_);
    or _11004_(_04544_, _04543_, _04538_);
    or _11005_(_04546_, _04544_, _04537_);
    or _11006_(_04547_, _04546_, _04522_);
    or _11007_(_04548_, _04478_, _04411_);
    and _11008_(_04549_, _04477_, _04437_);
    or _11009_(_04550_, _04432_, _03127_);
    and _11010_(_04551_, _04550_, _04470_);
    or _11011_(_04552_, _04551_, _04418_);
    and _11012_(_04553_, _04552_, _04463_);
    xnor _11013_(_04554_, _04553_, _04412_);
    or _11014_(_04555_, _04554_, _04549_);
    and _11015_(_04557_, _04555_, _04548_);
    xor _11016_(_04558_, _04557_, _00429_);
    or _11017_(_04559_, _04478_, _04417_);
    xnor _11018_(_04560_, _04551_, _04418_);
    or _11019_(_04561_, _04560_, _04549_);
    and _11020_(_04562_, _04561_, _04559_);
    xor _11021_(_04563_, _04562_, _00309_);
    or _11022_(_04564_, _04563_, _04558_);
    or _11023_(_04565_, _04478_, _04425_);
    or _11024_(_04566_, _04431_, _03127_);
    and _11025_(_04568_, _04566_, _04467_);
    xnor _11026_(_04569_, _04568_, _04426_);
    or _11027_(_04570_, _04569_, _04549_);
    and _11028_(_04571_, _04570_, _04565_);
    xor _11029_(_04572_, _04571_, _00183_);
    or _11030_(_04573_, _04478_, _04430_);
    xor _11031_(_04574_, _04431_, _03376_);
    or _11032_(_04575_, _04574_, _04549_);
    and _11033_(_04576_, _04575_, _04573_);
    xor _11034_(_04577_, _04576_, _06035_);
    or _11035_(_04579_, _04577_, _04572_);
    or _11036_(_04580_, _04579_, _04564_);
    not _11037_(_04581_, _04580_);
    xor _11038_(_04582_, _02984_, modulus[0]);
    and _11039_(_04583_, _04582_, _02985_);
    and _11040_(_04584_, _04583_, _02988_);
    nand _11041_(_04585_, _04584_, _04581_);
    nor _11042_(_04586_, _04585_, _04547_);
    nand _11043_(_04587_, _04586_, _05958_);
    or _11044_(_04588_, _04491_, modulus[12]);
    or _11045_(_04590_, _04542_, modulus[11]);
    or _11046_(_04591_, _04590_, _04538_);
    and _11047_(_04592_, _04591_, _04588_);
    or _11048_(_04593_, _04529_, modulus[10]);
    or _11049_(_04594_, _04535_, modulus[9]);
    or _11050_(_04595_, _04594_, _04530_);
    and _11051_(_04596_, _04595_, _04593_);
    or _11052_(_04597_, _04596_, _04544_);
    and _11053_(_04598_, _04597_, _04592_);
    or _11054_(_04599_, _04499_, modulus[8]);
    or _11055_(_04601_, _04505_, modulus[7]);
    or _11056_(_04602_, _04601_, _04500_);
    and _11057_(_04603_, _04602_, _04599_);
    or _11058_(_04604_, _04514_, modulus[6]);
    or _11059_(_04605_, _04519_, modulus[5]);
    or _11060_(_04606_, _04605_, _04515_);
    and _11061_(_04607_, _04606_, _04604_);
    or _11062_(_04608_, _04607_, _04507_);
    and _11063_(_04609_, _04608_, _04603_);
    or _11064_(_04610_, _04609_, _04546_);
    and _11065_(_04612_, _04610_, _04598_);
    or _11066_(_04613_, _04557_, modulus[4]);
    or _11067_(_04614_, _04562_, modulus[3]);
    or _11068_(_04615_, _04614_, _04558_);
    and _11069_(_04616_, _04615_, _04613_);
    or _11070_(_04617_, _04571_, modulus[2]);
    or _11071_(_04618_, _04576_, modulus[1]);
    or _11072_(_04619_, _04618_, _04572_);
    and _11073_(_04620_, _04619_, _04617_);
    or _11074_(_04621_, _04620_, _04564_);
    and _11075_(_04623_, _04621_, _04616_);
    and _11076_(_04624_, _02984_, modulus[0]);
    or _11077_(_04625_, _04624_, _04580_);
    and _11078_(_04626_, _04625_, _04623_);
    or _11079_(_04627_, _04626_, _04547_);
    nand _11080_(_04628_, _04627_, _04612_);
    and _11081_(_04629_, _04628_, _05957_);
    nand _11082_(_04630_, _04629_, _05956_);
    nand _11083_(_04631_, _04630_, _04587_);
    or _11084_(_04632_, _04631_, _04491_);
    or _11085_(_04634_, _04626_, _04522_);
    and _11086_(_04635_, _04634_, _04609_);
    or _11087_(_04636_, _04635_, _04537_);
    and _11088_(_04637_, _04636_, _04596_);
    or _11089_(_04638_, _04637_, _04543_);
    and _11090_(_04639_, _04638_, _04590_);
    xor _11091_(_04640_, _04639_, _04538_);
    nand _11092_(_04641_, _04640_, _04631_);
    and _11093_(_04642_, _04641_, _04632_);
    or _11094_(_04643_, _04631_, _04499_);
    or _11095_(_04645_, _04626_, _04521_);
    and _11096_(_04646_, _04645_, _04607_);
    or _11097_(_04647_, _04646_, _04506_);
    and _11098_(_04648_, _04647_, _04601_);
    xor _11099_(_04649_, _04648_, _04500_);
    nand _11100_(_04650_, _04649_, _04631_);
    and _11101_(_04651_, _04650_, _04643_);
    xor _11102_(_04652_, _04651_, _01048_);
    or _11103_(_04653_, _04631_, _04505_);
    and _11104_(_04654_, _04630_, _04587_);
    xnor _11105_(_04656_, _04646_, _04506_);
    or _11106_(_04657_, _04656_, _04654_);
    and _11107_(_04658_, _04657_, _04653_);
    xor _11108_(_04659_, _04658_, _00919_);
    or _11109_(_04660_, _04659_, _04652_);
    or _11110_(_04661_, _04631_, _04514_);
    or _11111_(_04662_, _04626_, _04520_);
    and _11112_(_04663_, _04662_, _04605_);
    xnor _11113_(_04664_, _04663_, _04515_);
    or _11114_(_04665_, _04664_, _04654_);
    and _11115_(_04667_, _04665_, _04661_);
    xor _11116_(_04668_, _04667_, _00797_);
    or _11117_(_04669_, _04631_, _04519_);
    xnor _11118_(_04670_, _04626_, _04520_);
    or _11119_(_04671_, _04670_, _04654_);
    and _11120_(_04672_, _04671_, _04669_);
    xor _11121_(_04673_, _04672_, _00673_);
    or _11122_(_04674_, _04673_, _04668_);
    or _11123_(_04675_, _04674_, _04660_);
    or _11124_(_04676_, _04631_, _04529_);
    or _11125_(_04678_, _04635_, _04536_);
    and _11126_(_04679_, _04678_, _04594_);
    xor _11127_(_04680_, _04679_, _04530_);
    nand _11128_(_04681_, _04680_, _04631_);
    and _11129_(_04682_, _04681_, _04676_);
    xor _11130_(_04683_, _04682_, _01328_);
    or _11131_(_04684_, _04631_, _04535_);
    xnor _11132_(_04685_, _04635_, _04536_);
    or _11133_(_04686_, _04685_, _04654_);
    and _11134_(_04687_, _04686_, _04684_);
    xor _11135_(_04689_, _04687_, _01181_);
    or _11136_(_04690_, _04689_, _04683_);
    xor _11137_(_04691_, _04642_, _01628_);
    or _11138_(_04692_, _04631_, _04542_);
    xor _11139_(_04693_, _04637_, _04543_);
    nand _11140_(_04694_, _04693_, _04631_);
    and _11141_(_04695_, _04694_, _04692_);
    xor _11142_(_04696_, _04695_, _01474_);
    or _11143_(_04697_, _04696_, _04691_);
    or _11144_(_04698_, _04697_, _04690_);
    nor _11145_(_04700_, _04698_, _04675_);
    or _11146_(_04701_, _04631_, _04557_);
    or _11147_(_04702_, _04624_, _04579_);
    and _11148_(_04703_, _04702_, _04620_);
    or _11149_(_04704_, _04703_, _04563_);
    and _11150_(_04705_, _04704_, _04614_);
    xnor _11151_(_04706_, _04705_, _04558_);
    or _11152_(_04707_, _04706_, _04654_);
    and _11153_(_04708_, _04707_, _04701_);
    xor _11154_(_04709_, _04708_, _00550_);
    or _11155_(_04711_, _04631_, _04562_);
    xnor _11156_(_04712_, _04703_, _04563_);
    or _11157_(_04713_, _04712_, _04654_);
    and _11158_(_04714_, _04713_, _04711_);
    xor _11159_(_04715_, _04714_, _00429_);
    or _11160_(_04716_, _04715_, _04709_);
    or _11161_(_04717_, _04631_, _04571_);
    or _11162_(_04718_, _04624_, _04577_);
    and _11163_(_04719_, _04718_, _04618_);
    xnor _11164_(_04720_, _04719_, _04572_);
    or _11165_(_04722_, _04720_, _04654_);
    and _11166_(_04723_, _04722_, _04717_);
    xor _11167_(_04724_, _04723_, _00309_);
    or _11168_(_04725_, _04631_, _04576_);
    xnor _11169_(_04726_, _04624_, _04577_);
    or _11170_(_04727_, _04726_, _04654_);
    and _11171_(_04728_, _04727_, _04725_);
    xor _11172_(_04729_, _04728_, _00183_);
    or _11173_(_04730_, _04729_, _04724_);
    or _11174_(_04731_, _04730_, _04716_);
    or _11175_(_04733_, _04631_, _02984_);
    or _11176_(_04734_, _04654_, _04582_);
    and _11177_(_04735_, _04734_, _04733_);
    xor _11178_(_04736_, _04735_, modulus[1]);
    xor _11179_(_04737_, _02985_, _05927_);
    not _11180_(_04738_, _04737_);
    and _11181_(_04739_, _04738_, _04736_);
    nand _11182_(_04740_, _04739_, _02988_);
    nor _11183_(_04741_, _04740_, _04731_);
    and _11184_(_04742_, _04741_, _04700_);
    nand _11185_(_04744_, _04742_, _06071_);
    or _11186_(_04745_, _04642_, modulus[13]);
    or _11187_(_04746_, _04695_, modulus[12]);
    or _11188_(_04747_, _04746_, _04691_);
    and _11189_(_04748_, _04747_, _04745_);
    or _11190_(_04749_, _04682_, modulus[11]);
    or _11191_(_04750_, _04687_, modulus[10]);
    or _11192_(_04751_, _04750_, _04683_);
    and _11193_(_04752_, _04751_, _04749_);
    or _11194_(_04753_, _04752_, _04697_);
    and _11195_(_04755_, _04753_, _04748_);
    or _11196_(_04756_, _04651_, modulus[9]);
    or _11197_(_04757_, _04658_, modulus[8]);
    or _11198_(_04758_, _04757_, _04652_);
    and _11199_(_04759_, _04758_, _04756_);
    or _11200_(_04760_, _04667_, modulus[7]);
    or _11201_(_04761_, _04672_, modulus[6]);
    or _11202_(_04762_, _04761_, _04668_);
    and _11203_(_04763_, _04762_, _04760_);
    or _11204_(_04764_, _04763_, _04660_);
    and _11205_(_04766_, _04764_, _04759_);
    or _11206_(_04767_, _04766_, _04698_);
    and _11207_(_04768_, _04767_, _04755_);
    or _11208_(_04769_, _04708_, modulus[5]);
    or _11209_(_04770_, _04714_, modulus[4]);
    or _11210_(_04771_, _04770_, _04709_);
    and _11211_(_04772_, _04771_, _04769_);
    or _11212_(_04773_, _04723_, modulus[3]);
    or _11213_(_04774_, _04728_, modulus[2]);
    or _11214_(_04775_, _04774_, _04724_);
    and _11215_(_04777_, _04775_, _04773_);
    or _11216_(_04778_, _04777_, _04716_);
    and _11217_(_04779_, _04778_, _04772_);
    or _11218_(_04780_, _04735_, modulus[1]);
    nor _11219_(_04781_, _02985_, modulus[0]);
    nand _11220_(_04782_, _04781_, _04736_);
    nand _11221_(_04783_, _04782_, _04780_);
    nor _11222_(_04784_, _04783_, _04739_);
    or _11223_(_04785_, _04784_, _04731_);
    nand _11224_(_04786_, _04785_, _04779_);
    nand _11225_(_04788_, _04786_, _04700_);
    nand _11226_(_04789_, _04788_, _04768_);
    nand _11227_(_04790_, _04789_, _06071_);
    nand _11228_(_04791_, _04790_, _04744_);
    or _11229_(_04792_, _04791_, _04642_);
    and _11230_(_04793_, _04790_, _04744_);
    and _11231_(_04794_, _04785_, _04779_);
    or _11232_(_04795_, _04794_, _04675_);
    and _11233_(_04796_, _04795_, _04766_);
    or _11234_(_04797_, _04796_, _04690_);
    and _11235_(_04799_, _04797_, _04752_);
    or _11236_(_04800_, _04799_, _04696_);
    nand _11237_(_04801_, _04800_, _04746_);
    xor _11238_(_04802_, _04801_, _04691_);
    or _11239_(_04803_, _04802_, _04793_);
    and _11240_(_04804_, _04803_, _04792_);
    or _11241_(_04805_, _04791_, _04651_);
    or _11242_(_04806_, _04794_, _04674_);
    and _11243_(_04807_, _04806_, _04763_);
    or _11244_(_04808_, _04807_, _04659_);
    nand _11245_(_04809_, _04808_, _04757_);
    xor _11246_(_04810_, _04809_, _04652_);
    or _11247_(_04811_, _04810_, _04793_);
    and _11248_(_04812_, _04811_, _04805_);
    xor _11249_(_04813_, _04812_, _01181_);
    or _11250_(_04814_, _04791_, _04658_);
    xnor _11251_(_04815_, _04807_, _04659_);
    or _11252_(_04816_, _04815_, _04793_);
    and _11253_(_04817_, _04816_, _04814_);
    xor _11254_(_04818_, _04817_, _01048_);
    or _11255_(_04820_, _04818_, _04813_);
    or _11256_(_04821_, _04791_, _04667_);
    or _11257_(_04822_, _04794_, _04673_);
    nand _11258_(_04823_, _04822_, _04761_);
    xor _11259_(_04824_, _04823_, _04668_);
    or _11260_(_04825_, _04824_, _04793_);
    and _11261_(_04826_, _04825_, _04821_);
    xor _11262_(_04827_, _04826_, _00919_);
    or _11263_(_04828_, _04791_, _04672_);
    xor _11264_(_04829_, _04786_, _04673_);
    or _11265_(_04831_, _04829_, _04793_);
    and _11266_(_04832_, _04831_, _04828_);
    xor _11267_(_04833_, _04832_, _00797_);
    or _11268_(_04834_, _04833_, _04827_);
    or _11269_(_04835_, _04834_, _04820_);
    or _11270_(_04836_, _04791_, _04682_);
    or _11271_(_04837_, _04796_, _04689_);
    nand _11272_(_04838_, _04837_, _04750_);
    xor _11273_(_04839_, _04838_, _04683_);
    or _11274_(_04840_, _04839_, _04793_);
    and _11275_(_04842_, _04840_, _04836_);
    xor _11276_(_04843_, _04842_, _01474_);
    or _11277_(_04844_, _04791_, _04687_);
    xnor _11278_(_04845_, _04796_, _04689_);
    or _11279_(_04846_, _04845_, _04793_);
    and _11280_(_04847_, _04846_, _04844_);
    xor _11281_(_04848_, _04847_, _01328_);
    or _11282_(_04849_, _04848_, _04843_);
    xor _11283_(_04850_, _04804_, _01789_);
    or _11284_(_04851_, _04791_, _04695_);
    xnor _11285_(_04853_, _04799_, _04696_);
    or _11286_(_04854_, _04853_, _04793_);
    and _11287_(_04855_, _04854_, _04851_);
    xor _11288_(_04856_, _04855_, _01628_);
    or _11289_(_04857_, _04856_, _04850_);
    or _11290_(_04858_, _04857_, _04849_);
    or _11291_(_04859_, _04858_, _04835_);
    or _11292_(_04860_, _04791_, _04708_);
    or _11293_(_04861_, _04784_, _04730_);
    and _11294_(_04862_, _04861_, _04777_);
    or _11295_(_04864_, _04862_, _04715_);
    nand _11296_(_04865_, _04864_, _04770_);
    xor _11297_(_04866_, _04865_, _04709_);
    or _11298_(_04867_, _04866_, _04793_);
    and _11299_(_04868_, _04867_, _04860_);
    xor _11300_(_04869_, _04868_, _00673_);
    or _11301_(_04870_, _04791_, _04714_);
    xnor _11302_(_04871_, _04862_, _04715_);
    or _11303_(_04872_, _04871_, _04793_);
    and _11304_(_04873_, _04872_, _04870_);
    xor _11305_(_04875_, _04873_, _00550_);
    or _11306_(_04876_, _04875_, _04869_);
    or _11307_(_04877_, _04791_, _04723_);
    or _11308_(_04878_, _04784_, _04729_);
    nand _11309_(_04879_, _04878_, _04774_);
    xor _11310_(_04880_, _04879_, _04724_);
    or _11311_(_04881_, _04880_, _04793_);
    and _11312_(_04882_, _04881_, _04877_);
    xor _11313_(_04883_, _04882_, _00429_);
    or _11314_(_04884_, _04791_, _04728_);
    xnor _11315_(_04886_, _04784_, _04729_);
    or _11316_(_04887_, _04886_, _04793_);
    and _11317_(_04888_, _04887_, _04884_);
    xor _11318_(_04889_, _04888_, _00309_);
    or _11319_(_04890_, _04889_, _04883_);
    nor _11320_(_04891_, _04890_, _04876_);
    or _11321_(_04892_, _04791_, _04735_);
    and _11322_(_04893_, _02985_, modulus[0]);
    xor _11323_(_04894_, _04893_, _04736_);
    or _11324_(_04895_, _04894_, _04793_);
    and _11325_(_04897_, _04895_, _04892_);
    xor _11326_(_04898_, _04897_, _00183_);
    or _11327_(_04899_, _04791_, _02985_);
    or _11328_(_04900_, _04793_, _04738_);
    and _11329_(_04901_, _04900_, _04899_);
    xor _11330_(_04902_, _04901_, _06035_);
    or _11331_(_04903_, _04902_, _04898_);
    xor _11332_(_04904_, _02987_, modulus[0]);
    nand _11333_(_04905_, _04904_, _02120_);
    nor _11334_(_04906_, _04905_, _04903_);
    nand _11335_(_04908_, _04906_, _04891_);
    nor _11336_(_04909_, _04908_, _04859_);
    or _11337_(_04910_, _04804_, modulus[14]);
    or _11338_(_04911_, _04855_, modulus[13]);
    or _11339_(_04912_, _04911_, _04850_);
    and _11340_(_04913_, _04912_, _04910_);
    or _11341_(_04914_, _04842_, modulus[12]);
    or _11342_(_04915_, _04847_, modulus[11]);
    or _11343_(_04916_, _04915_, _04843_);
    and _11344_(_04917_, _04916_, _04914_);
    or _11345_(_04919_, _04917_, _04857_);
    and _11346_(_04920_, _04919_, _04913_);
    or _11347_(_04921_, _04812_, modulus[10]);
    or _11348_(_04922_, _04817_, modulus[9]);
    or _11349_(_04923_, _04922_, _04813_);
    and _11350_(_04924_, _04923_, _04921_);
    or _11351_(_04925_, _04826_, modulus[8]);
    or _11352_(_04926_, _04832_, modulus[7]);
    or _11353_(_04927_, _04926_, _04827_);
    and _11354_(_04928_, _04927_, _04925_);
    or _11355_(_04930_, _04928_, _04820_);
    and _11356_(_04931_, _04930_, _04924_);
    or _11357_(_04932_, _04931_, _04858_);
    and _11358_(_04933_, _04932_, _04920_);
    or _11359_(_04934_, _04868_, modulus[6]);
    or _11360_(_04935_, _04873_, modulus[5]);
    or _11361_(_04936_, _04935_, _04869_);
    and _11362_(_04937_, _04936_, _04934_);
    or _11363_(_04938_, _04882_, modulus[4]);
    or _11364_(_04939_, _04888_, modulus[3]);
    or _11365_(_04941_, _04939_, _04883_);
    and _11366_(_04942_, _04941_, _04938_);
    or _11367_(_04943_, _04942_, _04876_);
    and _11368_(_04944_, _04943_, _04937_);
    not _11369_(_04945_, _04891_);
    or _11370_(_04946_, _04897_, modulus[2]);
    or _11371_(_04947_, _04901_, modulus[1]);
    or _11372_(_04948_, _04947_, _04898_);
    and _11373_(_04949_, _04948_, _04946_);
    and _11374_(_04950_, _02987_, modulus[0]);
    or _11375_(_04952_, _04950_, _04903_);
    and _11376_(_04953_, _04952_, _04949_);
    or _11377_(_04954_, _04953_, _04945_);
    and _11378_(_04955_, _04954_, _04944_);
    or _11379_(_04956_, _04955_, _04859_);
    and _11380_(_04957_, _04956_, _04933_);
    or _11381_(_04958_, _04955_, _04835_);
    and _11382_(_04959_, _04958_, _04931_);
    or _11383_(_04960_, _04959_, _04849_);
    and _11384_(_04961_, _04960_, _04917_);
    or _11385_(_04963_, _04961_, _04856_);
    nand _11386_(_04964_, _04963_, _04911_);
    xor _11387_(_04965_, _04964_, _04850_);
    and _11388_(_04966_, _04804_, modulus[15]);
    nand _11389_(_04967_, _04909_, _05956_);
    or _11390_(_04968_, _04957_, modulus[15]);
    nand _11391_(_04969_, _04968_, _04967_);
    or _11392_(_04970_, _04969_, _04804_);
    and _11393_(_04971_, _04968_, _04967_);
    or _11394_(_04972_, _04965_, _04971_);
    and _11395_(_04974_, _04972_, _04970_);
    xor _11396_(_04975_, _04974_, _05956_);
    or _11397_(_04976_, _04969_, _04855_);
    xnor _11398_(_04977_, _04961_, _04856_);
    or _11399_(_04978_, _04977_, _04971_);
    and _11400_(_04979_, _04978_, _04976_);
    nand _11401_(_04980_, _04979_, modulus[14]);
    nor _11402_(_04981_, _04980_, _04975_);
    nor _11403_(_04982_, _04981_, _04966_);
    xor _11404_(_04983_, _04979_, _01789_);
    nor _11405_(_04985_, _04983_, _04975_);
    not _11406_(_04986_, _04985_);
    or _11407_(_04987_, _04969_, _04842_);
    or _11408_(_04988_, _04959_, _04848_);
    nand _11409_(_04989_, _04988_, _04915_);
    xor _11410_(_04990_, _04989_, _04843_);
    or _11411_(_04991_, _04990_, _04971_);
    and _11412_(_04992_, _04991_, _04987_);
    and _11413_(_04993_, _04992_, modulus[13]);
    xor _11414_(_04994_, _04992_, _01628_);
    not _11415_(_04996_, _04994_);
    or _11416_(_04997_, _04969_, _04847_);
    xnor _11417_(_04998_, _04959_, _04848_);
    or _11418_(_04999_, _04998_, _04971_);
    and _11419_(_05000_, _04999_, _04997_);
    and _11420_(_05001_, _05000_, modulus[12]);
    and _11421_(_05002_, _05001_, _04996_);
    nor _11422_(_05003_, _05002_, _04993_);
    or _11423_(_05004_, _05003_, _04986_);
    and _11424_(_05005_, _05004_, _04982_);
    xor _11425_(_05007_, _05000_, _01474_);
    nor _11426_(_05008_, _05007_, _04994_);
    and _11427_(_05009_, _05008_, _04985_);
    or _11428_(_05010_, _04969_, _04812_);
    or _11429_(_05011_, _04955_, _04834_);
    and _11430_(_05012_, _05011_, _04928_);
    or _11431_(_05013_, _05012_, _04818_);
    nand _11432_(_05014_, _05013_, _04922_);
    xor _11433_(_05015_, _05014_, _04813_);
    or _11434_(_05016_, _05015_, _04971_);
    and _11435_(_05018_, _05016_, _05010_);
    and _11436_(_05019_, _05018_, modulus[11]);
    xor _11437_(_05020_, _05018_, _01328_);
    or _11438_(_05021_, _04969_, _04817_);
    xnor _11439_(_05022_, _05012_, _04818_);
    or _11440_(_05023_, _05022_, _04971_);
    and _11441_(_05024_, _05023_, _05021_);
    nand _11442_(_05025_, _05024_, modulus[10]);
    nor _11443_(_05026_, _05025_, _05020_);
    nor _11444_(_05027_, _05026_, _05019_);
    not _11445_(_05029_, _05027_);
    xor _11446_(_05030_, _05024_, _01181_);
    or _11447_(_05031_, _05030_, _05020_);
    or _11448_(_05032_, _04969_, _04826_);
    or _11449_(_05033_, _04955_, _04833_);
    nand _11450_(_05034_, _05033_, _04926_);
    xor _11451_(_05035_, _05034_, _04827_);
    or _11452_(_05036_, _05035_, _04971_);
    and _11453_(_05037_, _05036_, _05032_);
    nand _11454_(_05038_, _05037_, modulus[9]);
    xor _11455_(_05040_, _05037_, _01048_);
    or _11456_(_05041_, _04969_, _04832_);
    xnor _11457_(_05042_, _04955_, _04833_);
    or _11458_(_05043_, _05042_, _04971_);
    and _11459_(_05044_, _05043_, _05041_);
    nand _11460_(_05045_, _05044_, modulus[8]);
    or _11461_(_05046_, _05045_, _05040_);
    and _11462_(_05047_, _05046_, _05038_);
    nor _11463_(_05048_, _05047_, _05031_);
    or _11464_(_05049_, _05048_, _05029_);
    nand _11465_(_05051_, _05049_, _05009_);
    and _11466_(_05052_, _05051_, _05005_);
    xor _11467_(_05053_, _05044_, _00919_);
    or _11468_(_05054_, _05053_, _05040_);
    or _11469_(_05055_, _05054_, _05031_);
    not _11470_(_05056_, _05055_);
    and _11471_(_05057_, _05056_, _05009_);
    or _11472_(_05058_, _04969_, _04868_);
    or _11473_(_05059_, _04953_, _04890_);
    and _11474_(_05060_, _05059_, _04942_);
    or _11475_(_05062_, _05060_, _04875_);
    nand _11476_(_05063_, _05062_, _04935_);
    xor _11477_(_05064_, _05063_, _04869_);
    or _11478_(_05065_, _05064_, _04971_);
    and _11479_(_05066_, _05065_, _05058_);
    and _11480_(_05067_, _05066_, modulus[7]);
    xor _11481_(_05068_, _05066_, _00797_);
    or _11482_(_05069_, _04969_, _04873_);
    xnor _11483_(_05070_, _05060_, _04875_);
    or _11484_(_05071_, _05070_, _04971_);
    and _11485_(_05073_, _05071_, _05069_);
    nand _11486_(_05074_, _05073_, modulus[6]);
    nor _11487_(_05075_, _05074_, _05068_);
    nor _11488_(_05076_, _05075_, _05067_);
    not _11489_(_05077_, _05076_);
    xor _11490_(_05078_, _05073_, _00673_);
    or _11491_(_05079_, _05078_, _05068_);
    or _11492_(_05080_, _04969_, _04882_);
    or _11493_(_05081_, _04953_, _04889_);
    nand _11494_(_05082_, _05081_, _04939_);
    xor _11495_(_05084_, _05082_, _04883_);
    or _11496_(_05085_, _05084_, _04971_);
    and _11497_(_05086_, _05085_, _05080_);
    nand _11498_(_05087_, _05086_, modulus[5]);
    xor _11499_(_05088_, _05086_, _00550_);
    or _11500_(_05089_, _04969_, _04888_);
    xnor _11501_(_05090_, _04953_, _04889_);
    or _11502_(_05091_, _05090_, _04971_);
    and _11503_(_05092_, _05091_, _05089_);
    nand _11504_(_05093_, _05092_, modulus[4]);
    or _11505_(_05095_, _05093_, _05088_);
    and _11506_(_05096_, _05095_, _05087_);
    nor _11507_(_05097_, _05096_, _05079_);
    nor _11508_(_05098_, _05097_, _05077_);
    xor _11509_(_05099_, _05092_, _00429_);
    or _11510_(_05100_, _05099_, _05088_);
    or _11511_(_05101_, _05100_, _05079_);
    or _11512_(_05102_, _04969_, _04897_);
    or _11513_(_05103_, _04950_, _04902_);
    nand _11514_(_05104_, _05103_, _04947_);
    xor _11515_(_05106_, _05104_, _04898_);
    or _11516_(_05107_, _05106_, _04971_);
    and _11517_(_05108_, _05107_, _05102_);
    nand _11518_(_05109_, _05108_, modulus[3]);
    xor _11519_(_05110_, _05108_, _00309_);
    or _11520_(_05111_, _04969_, _04901_);
    xnor _11521_(_05112_, _04950_, _04902_);
    or _11522_(_05113_, _05112_, _04971_);
    and _11523_(_05114_, _05113_, _05111_);
    nand _11524_(_05115_, _05114_, modulus[2]);
    or _11525_(_05117_, _05115_, _05110_);
    and _11526_(_05118_, _05117_, _05109_);
    xor _11527_(_05119_, _05114_, _00183_);
    or _11528_(_05120_, _05119_, _05110_);
    or _11529_(_05121_, _04969_, _02987_);
    or _11530_(_05122_, _04971_, _04904_);
    and _11531_(_05123_, _05122_, _05121_);
    nand _11532_(_05124_, _05123_, modulus[1]);
    xor _11533_(_05125_, _05123_, _06035_);
    and _11534_(_05126_, _02119_, _05927_);
    or _11535_(_05128_, _05126_, _05125_);
    and _11536_(_05129_, _05128_, _05124_);
    or _11537_(_05130_, _05129_, _05120_);
    and _11538_(_05131_, _05130_, _05118_);
    or _11539_(_05132_, _05131_, _05101_);
    nand _11540_(_05133_, _05132_, _05098_);
    nand _11541_(_05134_, _05133_, _05057_);
    and _11542_(_05135_, _05134_, _05052_);
    not _11543_(_05136_, _05101_);
    not _11544_(_05137_, _05120_);
    xor _11545_(_05139_, _02119_, modulus[0]);
    nor _11546_(_05140_, _05139_, _05125_);
    and _11547_(_05141_, _05140_, _05137_);
    and _11548_(_05142_, _05141_, _05136_);
    and _11549_(_05143_, _05142_, _05057_);
    or _11550_(_05144_, _05143_, _05135_);
    nor _11551_(_05145_, _05144_, _02120_);
    and _11552_(_05146_, _05144_, _05139_);
    or _11553_(_05147_, _05146_, _05145_);
    and _11554_(_05148_, _05147_, exp_counter[0]);
    and _11555_(_05150_, _05148_, _02084_);
    and _11556_(_05151_, _05150_, rsa_active);
    or _11557_(_05152_, _05151_, _01160_);
    and _11558_(_05153_, _05152_, _02116_);
    or _11559_(_00057_, _05153_, _02118_);
    and _11560_(_05154_, _02117_, accumulator[1]);
    nor _11561_(_05155_, _05144_, _05123_);
    nor _11562_(_05156_, _02119_, _05927_);
    xor _11563_(_05157_, _05156_, _05125_);
    and _11564_(_05158_, _05157_, _05144_);
    or _11565_(_05160_, _05158_, _05155_);
    and _11566_(_05161_, _05160_, exp_counter[0]);
    and _11567_(_05162_, _05161_, _02084_);
    and _11568_(_05163_, _05162_, rsa_active);
    and _11569_(_05164_, _05163_, _02093_);
    and _11570_(_05165_, _05164_, _02116_);
    or _11571_(_00058_, _05165_, _05154_);
    and _11572_(_05166_, _02117_, accumulator[2]);
    nor _11573_(_05167_, _05144_, _05114_);
    or _11574_(_05168_, _05123_, modulus[1]);
    or _11575_(_05170_, _05156_, _05125_);
    and _11576_(_05171_, _05170_, _05168_);
    xor _11577_(_05172_, _05171_, _05119_);
    and _11578_(_05173_, _05172_, _05144_);
    or _11579_(_05174_, _05173_, _05167_);
    and _11580_(_05175_, _05174_, exp_counter[0]);
    and _11581_(_05176_, _05175_, _02084_);
    and _11582_(_05177_, _05176_, rsa_active);
    and _11583_(_05178_, _05177_, _02093_);
    and _11584_(_05179_, _05178_, _02116_);
    or _11585_(_00059_, _05179_, _05166_);
    and _11586_(_05181_, _02117_, accumulator[3]);
    nor _11587_(_05182_, _05144_, _05108_);
    or _11588_(_05183_, _05114_, modulus[2]);
    or _11589_(_05184_, _05171_, _05119_);
    and _11590_(_05185_, _05184_, _05183_);
    xor _11591_(_05186_, _05185_, _05110_);
    and _11592_(_05187_, _05186_, _05144_);
    or _11593_(_05188_, _05187_, _05182_);
    and _11594_(_05189_, _05188_, exp_counter[0]);
    and _11595_(_05191_, _05189_, _02084_);
    and _11596_(_05192_, _05191_, rsa_active);
    and _11597_(_05193_, _05192_, _02093_);
    and _11598_(_05194_, _05193_, _02116_);
    or _11599_(_00060_, _05194_, _05181_);
    and _11600_(_05195_, _02117_, accumulator[4]);
    nor _11601_(_05196_, _05144_, _05092_);
    or _11602_(_05197_, _05108_, modulus[3]);
    or _11603_(_05198_, _05183_, _05110_);
    and _11604_(_05199_, _05198_, _05197_);
    or _11605_(_05201_, _05171_, _05120_);
    and _11606_(_05202_, _05201_, _05199_);
    xor _11607_(_05203_, _05202_, _05099_);
    and _11608_(_05204_, _05203_, _05144_);
    or _11609_(_05205_, _05204_, _05196_);
    and _11610_(_05206_, _05205_, exp_counter[0]);
    and _11611_(_05207_, _05206_, _02084_);
    and _11612_(_05208_, _05207_, rsa_active);
    and _11613_(_05209_, _05208_, _02093_);
    and _11614_(_05210_, _05209_, _02116_);
    or _11615_(_00061_, _05210_, _05195_);
    and _11616_(_05212_, _02117_, accumulator[5]);
    nor _11617_(_05213_, _05144_, _05086_);
    or _11618_(_05214_, _05092_, modulus[4]);
    or _11619_(_05215_, _05202_, _05099_);
    and _11620_(_05216_, _05215_, _05214_);
    xor _11621_(_05217_, _05216_, _05088_);
    and _11622_(_05218_, _05217_, _05144_);
    or _11623_(_05219_, _05218_, _05213_);
    and _11624_(_05220_, _05219_, exp_counter[0]);
    and _11625_(_05222_, _05220_, _02084_);
    and _11626_(_05223_, _05222_, rsa_active);
    and _11627_(_05224_, _05223_, _02093_);
    and _11628_(_05225_, _05224_, _02116_);
    or _11629_(_00062_, _05225_, _05212_);
    and _11630_(_05226_, _02117_, accumulator[6]);
    nor _11631_(_05227_, _05144_, _05073_);
    or _11632_(_05228_, _05086_, modulus[5]);
    or _11633_(_05229_, _05214_, _05088_);
    and _11634_(_05230_, _05229_, _05228_);
    or _11635_(_05232_, _05202_, _05100_);
    and _11636_(_05233_, _05232_, _05230_);
    xor _11637_(_05234_, _05233_, _05078_);
    and _11638_(_05235_, _05234_, _05144_);
    or _11639_(_05236_, _05235_, _05227_);
    and _11640_(_05237_, _05236_, exp_counter[0]);
    and _11641_(_05238_, _05237_, _02084_);
    and _11642_(_05239_, _05238_, rsa_active);
    and _11643_(_05240_, _05239_, _02093_);
    and _11644_(_05241_, _05240_, _02116_);
    or _11645_(_00063_, _05241_, _05226_);
    and _11646_(_05243_, _02117_, accumulator[7]);
    nor _11647_(_05244_, _05144_, _05066_);
    or _11648_(_05245_, _05073_, modulus[6]);
    or _11649_(_05246_, _05233_, _05078_);
    and _11650_(_05247_, _05246_, _05245_);
    xor _11651_(_05248_, _05247_, _05068_);
    and _11652_(_05249_, _05248_, _05144_);
    or _11653_(_05250_, _05249_, _05244_);
    and _11654_(_05251_, _05250_, exp_counter[0]);
    and _11655_(_05253_, _05251_, _02084_);
    and _11656_(_05254_, _05253_, rsa_active);
    and _11657_(_05255_, _05254_, _02093_);
    and _11658_(_05256_, _05255_, _02116_);
    or _11659_(_00064_, _05256_, _05243_);
    and _11660_(_05257_, _02117_, accumulator[8]);
    nor _11661_(_05258_, _05144_, _05044_);
    or _11662_(_05259_, _05066_, modulus[7]);
    or _11663_(_05260_, _05245_, _05068_);
    and _11664_(_05261_, _05260_, _05259_);
    or _11665_(_05263_, _05230_, _05079_);
    and _11666_(_05264_, _05263_, _05261_);
    or _11667_(_05265_, _05202_, _05101_);
    and _11668_(_05266_, _05265_, _05264_);
    xor _11669_(_05267_, _05266_, _05053_);
    and _11670_(_05268_, _05267_, _05144_);
    or _11671_(_05269_, _05268_, _05258_);
    and _11672_(_05270_, _05269_, exp_counter[0]);
    and _11673_(_05271_, _05270_, _02084_);
    and _11674_(_05272_, _05271_, rsa_active);
    and _11675_(_05274_, _05272_, _02093_);
    and _11676_(_05275_, _05274_, _02116_);
    or _11677_(_00065_, _05275_, _05257_);
    and _11678_(_05276_, _02117_, accumulator[9]);
    nor _11679_(_05277_, _05144_, _05037_);
    or _11680_(_05278_, _05044_, modulus[8]);
    or _11681_(_05279_, _05266_, _05053_);
    and _11682_(_05280_, _05279_, _05278_);
    xor _11683_(_05281_, _05280_, _05040_);
    and _11684_(_05282_, _05281_, _05144_);
    or _11685_(_05284_, _05282_, _05277_);
    and _11686_(_05285_, _05284_, exp_counter[0]);
    and _11687_(_05286_, _05285_, _02084_);
    and _11688_(_05287_, _05286_, rsa_active);
    and _11689_(_05288_, _05287_, _02093_);
    and _11690_(_05289_, _05288_, _02116_);
    or _11691_(_00066_, _05289_, _05276_);
    and _11692_(_05290_, _02117_, accumulator[10]);
    nor _11693_(_05291_, _05144_, _05024_);
    or _11694_(_05292_, _05037_, modulus[9]);
    or _11695_(_05294_, _05278_, _05040_);
    and _11696_(_05295_, _05294_, _05292_);
    or _11697_(_05296_, _05266_, _05054_);
    and _11698_(_05297_, _05296_, _05295_);
    xor _11699_(_05298_, _05297_, _05030_);
    and _11700_(_05299_, _05298_, _05144_);
    or _11701_(_05300_, _05299_, _05291_);
    and _11702_(_05301_, _05300_, exp_counter[0]);
    and _11703_(_05302_, _05301_, _02084_);
    and _11704_(_05303_, _05302_, rsa_active);
    and _11705_(_05305_, _05303_, _02093_);
    and _11706_(_05306_, _05305_, _02116_);
    or _11707_(_00067_, _05306_, _05290_);
    and _11708_(_05307_, _02117_, accumulator[11]);
    nor _11709_(_05308_, _05144_, _05018_);
    or _11710_(_05309_, _05024_, modulus[10]);
    or _11711_(_05310_, _05297_, _05030_);
    and _11712_(_05311_, _05310_, _05309_);
    xor _11713_(_05312_, _05311_, _05020_);
    and _11714_(_05313_, _05312_, _05144_);
    or _11715_(_05315_, _05313_, _05308_);
    and _11716_(_05316_, _05315_, exp_counter[0]);
    and _11717_(_05317_, _05316_, _02084_);
    and _11718_(_05318_, _05317_, rsa_active);
    and _11719_(_05319_, _05318_, _02093_);
    and _11720_(_05320_, _05319_, _02116_);
    or _11721_(_00068_, _05320_, _05307_);
    and _11722_(_05321_, _02117_, accumulator[12]);
    nor _11723_(_05322_, _05144_, _05000_);
    or _11724_(_05323_, _05018_, modulus[11]);
    or _11725_(_05325_, _05309_, _05020_);
    and _11726_(_05326_, _05325_, _05323_);
    or _11727_(_05327_, _05295_, _05031_);
    and _11728_(_05328_, _05327_, _05326_);
    or _11729_(_05329_, _05266_, _05055_);
    and _11730_(_05330_, _05329_, _05328_);
    xor _11731_(_05331_, _05330_, _05007_);
    and _11732_(_05332_, _05331_, _05144_);
    or _11733_(_05333_, _05332_, _05322_);
    and _11734_(_05334_, _05333_, exp_counter[0]);
    and _11735_(_05336_, _05334_, _02084_);
    and _11736_(_05337_, _05336_, rsa_active);
    and _11737_(_05338_, _05337_, _02093_);
    and _11738_(_05339_, _05338_, _02116_);
    or _11739_(_00069_, _05339_, _05321_);
    and _11740_(_05340_, _02117_, accumulator[13]);
    nor _11741_(_05341_, _05144_, _04992_);
    or _11742_(_05342_, _05000_, modulus[12]);
    or _11743_(_05343_, _05330_, _05007_);
    and _11744_(_05344_, _05343_, _05342_);
    xor _11745_(_05346_, _05344_, _04994_);
    and _11746_(_05347_, _05346_, _05144_);
    or _11747_(_05348_, _05347_, _05341_);
    and _11748_(_05349_, _05348_, exp_counter[0]);
    and _11749_(_05350_, _05349_, _02084_);
    and _11750_(_05351_, _05350_, rsa_active);
    and _11751_(_05352_, _05351_, _02093_);
    and _11752_(_05353_, _05352_, _02116_);
    or _11753_(_00070_, _05353_, _05340_);
    and _11754_(_05354_, _02117_, accumulator[14]);
    nor _11755_(_05356_, _05144_, _04979_);
    or _11756_(_05357_, _04992_, modulus[13]);
    or _11757_(_05358_, _05342_, _04994_);
    and _11758_(_05359_, _05358_, _05357_);
    not _11759_(_05360_, _05008_);
    or _11760_(_05361_, _05330_, _05360_);
    and _11761_(_05362_, _05361_, _05359_);
    xor _11762_(_05363_, _05362_, _04983_);
    and _11763_(_05364_, _05363_, _05144_);
    or _11764_(_05365_, _05364_, _05356_);
    and _11765_(_05367_, _05365_, exp_counter[0]);
    and _11766_(_05368_, _05367_, _02084_);
    and _11767_(_05369_, _05368_, rsa_active);
    and _11768_(_05370_, _05369_, _02093_);
    and _11769_(_05371_, _05370_, _02116_);
    or _11770_(_00071_, _05371_, _05354_);
    and _11771_(_05372_, _02117_, accumulator[15]);
    nor _11772_(_05373_, _05144_, _04974_);
    or _11773_(_05374_, _04979_, modulus[14]);
    or _11774_(_05375_, _05362_, _04983_);
    and _11775_(_05377_, _05375_, _05374_);
    xor _11776_(_05378_, _05377_, _04975_);
    and _11777_(_05379_, _05378_, _05144_);
    or _11778_(_05380_, _05379_, _05373_);
    and _11779_(_05381_, _05380_, exp_counter[0]);
    and _11780_(_05382_, _05381_, _02084_);
    and _11781_(_05383_, _05382_, rsa_active);
    and _11782_(_05384_, _05383_, _02093_);
    and _11783_(_05385_, _05384_, _02116_);
    or _11784_(_00072_, _05385_, _05372_);
    nor _11785_(_05387_, _02089_, _05865_);
    and _11786_(_05388_, _02079_, _02057_);
    and _11787_(_05389_, modulus[0], _01138_);
    xnor _11788_(_05390_, _05389_, _02059_);
    nor _11789_(_05391_, _05390_, _02079_);
    or _11790_(_05392_, _05391_, _05388_);
    and _11791_(_05393_, _05392_, _02084_);
    and _11792_(_05394_, _05393_, rsa_active);
    and _11793_(_05395_, _05394_, _02093_);
    and _11794_(_05396_, _01160_, message[1]);
    or _11795_(_05398_, _05396_, _05395_);
    and _11796_(_05399_, _05398_, _02089_);
    or _11797_(_00073_, _05399_, _05387_);
    nor _11798_(_05400_, _02089_, _05806_);
    nor _11799_(_05401_, _02095_, _02051_);
    nand _11800_(_05402_, _02057_, _06035_);
    or _11801_(_05403_, _05389_, _02059_);
    and _11802_(_05404_, _05403_, _05402_);
    xnor _11803_(_05405_, _05404_, _02055_);
    nor _11804_(_05406_, _05405_, _02079_);
    or _11805_(_05408_, _05406_, _05401_);
    and _11806_(_05409_, _05408_, _02084_);
    and _11807_(_05410_, _05409_, rsa_active);
    and _11808_(_05411_, _05410_, _02093_);
    and _11809_(_05412_, _01160_, message[2]);
    or _11810_(_05413_, _05412_, _05411_);
    and _11811_(_05414_, _05413_, _02089_);
    or _11812_(_00074_, _05414_, _05400_);
    nor _11813_(_05415_, _02089_, _05773_);
    nor _11814_(_05416_, _02095_, _02044_);
    or _11815_(_05418_, _02051_, modulus[2]);
    or _11816_(_05419_, _05404_, _02055_);
    and _11817_(_05420_, _05419_, _05418_);
    xnor _11818_(_05421_, _05420_, _02046_);
    nor _11819_(_05422_, _05421_, _02079_);
    or _11820_(_05423_, _05422_, _05416_);
    and _11821_(_05424_, _05423_, _02084_);
    and _11822_(_05425_, _05424_, rsa_active);
    and _11823_(_05426_, _05425_, _02093_);
    and _11824_(_05427_, _01160_, message[3]);
    or _11825_(_05429_, _05427_, _05426_);
    and _11826_(_05430_, _05429_, _02089_);
    or _11827_(_00075_, _05430_, _05415_);
    nor _11828_(_05431_, _02089_, _05417_);
    nor _11829_(_05432_, _02095_, _02027_);
    or _11830_(_05433_, _02044_, modulus[3]);
    or _11831_(_05434_, _05418_, _02046_);
    and _11832_(_05435_, _05434_, _05433_);
    or _11833_(_05436_, _05404_, _02056_);
    and _11834_(_05437_, _05436_, _05435_);
    xnor _11835_(_05439_, _05437_, _02035_);
    nor _11836_(_05440_, _05439_, _02079_);
    or _11837_(_05441_, _05440_, _05432_);
    and _11838_(_05442_, _05441_, _02084_);
    and _11839_(_05443_, _05442_, rsa_active);
    and _11840_(_05444_, _05443_, _02093_);
    and _11841_(_05445_, _01160_, message[4]);
    or _11842_(_05446_, _05445_, _05444_);
    and _11843_(_05447_, _05446_, _02089_);
    or _11844_(_00076_, _05447_, _05431_);
    nor _11845_(_05449_, _02089_, _04215_);
    nor _11846_(_05450_, _02095_, _02021_);
    or _11847_(_05451_, _02027_, modulus[4]);
    or _11848_(_05452_, _05437_, _02035_);
    and _11849_(_05453_, _05452_, _05451_);
    xnor _11850_(_05454_, _05453_, _02023_);
    nor _11851_(_05455_, _05454_, _02079_);
    or _11852_(_05456_, _05455_, _05450_);
    and _11853_(_05457_, _05456_, _02084_);
    and _11854_(_05458_, _05457_, rsa_active);
    and _11855_(_05460_, _05458_, _02093_);
    and _11856_(_05461_, _01160_, message[5]);
    or _11857_(_05462_, _05461_, _05460_);
    and _11858_(_05463_, _05462_, _02089_);
    or _11859_(_00077_, _05463_, _05449_);
    and _11860_(_05464_, _02090_, base[6]);
    nor _11861_(_05465_, _02095_, _02009_);
    or _11862_(_05466_, _02021_, modulus[5]);
    or _11863_(_05467_, _05451_, _02023_);
    and _11864_(_05468_, _05467_, _05466_);
    or _11865_(_05470_, _05437_, _02036_);
    and _11866_(_05471_, _05470_, _05468_);
    xnor _11867_(_05472_, _05471_, _02013_);
    nor _11868_(_05473_, _05472_, _02079_);
    or _11869_(_05474_, _05473_, _05465_);
    and _11870_(_05475_, _05474_, _02084_);
    and _11871_(_05476_, _05475_, rsa_active);
    and _11872_(_05477_, _05476_, _02093_);
    and _11873_(_05478_, _01160_, message[6]);
    or _11874_(_05479_, _05478_, _05477_);
    and _11875_(_05481_, _05479_, _02089_);
    or _11876_(_00078_, _05481_, _05464_);
    nor _11877_(_05482_, _02089_, _01731_);
    nor _11878_(_05483_, _02095_, _02002_);
    or _11879_(_05484_, _02009_, modulus[6]);
    or _11880_(_05485_, _05471_, _02013_);
    and _11881_(_05486_, _05485_, _05484_);
    xnor _11882_(_05487_, _05486_, _02004_);
    nor _11883_(_05488_, _05487_, _02079_);
    or _11884_(_05489_, _05488_, _05483_);
    and _11885_(_05491_, _05489_, _02084_);
    and _11886_(_05492_, _05491_, rsa_active);
    and _11887_(_05493_, _05492_, _02093_);
    and _11888_(_05494_, _01160_, message[7]);
    or _11889_(_05495_, _05494_, _05493_);
    and _11890_(_05496_, _05495_, _02089_);
    or _11891_(_00079_, _05496_, _05482_);
    and _11892_(_05497_, _02090_, base[8]);
    nor _11893_(_05498_, _02095_, _01979_);
    or _11894_(_05499_, _02002_, modulus[7]);
    or _11895_(_05501_, _05484_, _02004_);
    and _11896_(_05502_, _05501_, _05499_);
    or _11897_(_05503_, _05468_, _02014_);
    and _11898_(_05504_, _05503_, _05502_);
    or _11899_(_05505_, _05437_, _02037_);
    and _11900_(_05506_, _05505_, _05504_);
    xnor _11901_(_05507_, _05506_, _01989_);
    nor _11902_(_05508_, _05507_, _02079_);
    or _11903_(_05509_, _05508_, _05498_);
    and _11904_(_05510_, _05509_, _02084_);
    and _11905_(_05512_, _05510_, rsa_active);
    and _11906_(_05513_, _05512_, _02093_);
    and _11907_(_05514_, _01160_, message[8]);
    or _11908_(_05515_, _05514_, _05513_);
    and _11909_(_05516_, _05515_, _02089_);
    or _11910_(_00080_, _05516_, _05497_);
    and _11911_(_05517_, _02090_, base[9]);
    nor _11912_(_05518_, _02095_, _01972_);
    or _11913_(_05519_, _01979_, modulus[8]);
    or _11914_(_05520_, _05506_, _01989_);
    and _11915_(_05522_, _05520_, _05519_);
    xnor _11916_(_05523_, _05522_, _01975_);
    nor _11917_(_05524_, _05523_, _02079_);
    or _11918_(_05525_, _05524_, _05518_);
    and _11919_(_05526_, _05525_, _02084_);
    and _11920_(_05527_, _05526_, rsa_active);
    and _11921_(_05528_, _05527_, _02093_);
    and _11922_(_05529_, _01160_, message[9]);
    or _11923_(_05530_, _05529_, _05528_);
    and _11924_(_05531_, _05530_, _02089_);
    or _11925_(_00081_, _05531_, _05517_);
    and _11926_(_05533_, _02090_, base[10]);
    nor _11927_(_05534_, _02095_, _01960_);
    or _11928_(_05535_, _01972_, modulus[9]);
    or _11929_(_05536_, _05519_, _01975_);
    and _11930_(_05537_, _05536_, _05535_);
    or _11931_(_05538_, _05506_, _01990_);
    and _11932_(_05539_, _05538_, _05537_);
    xnor _11933_(_05540_, _05539_, _01965_);
    nor _11934_(_05541_, _05540_, _02079_);
    or _11935_(_05543_, _05541_, _05534_);
    and _11936_(_05544_, _05543_, _02084_);
    and _11937_(_05545_, _05544_, rsa_active);
    and _11938_(_05546_, _05545_, _02093_);
    and _11939_(_05547_, _01160_, message[10]);
    or _11940_(_05548_, _05547_, _05546_);
    and _11941_(_05549_, _05548_, _02089_);
    or _11942_(_00082_, _05549_, _05533_);
    and _11943_(_05550_, _02090_, base[11]);
    nor _11944_(_05551_, _02095_, _01954_);
    or _11945_(_05553_, _01960_, modulus[10]);
    or _11946_(_05554_, _05539_, _01965_);
    and _11947_(_05555_, _05554_, _05553_);
    xnor _11948_(_05556_, _05555_, _01956_);
    nor _11949_(_05557_, _05556_, _02079_);
    or _11950_(_05558_, _05557_, _05551_);
    and _11951_(_05559_, _05558_, _02084_);
    and _11952_(_05560_, _05559_, rsa_active);
    and _11953_(_05561_, _05560_, _02093_);
    and _11954_(_05562_, _01160_, message[11]);
    or _11955_(_05564_, _05562_, _05561_);
    and _11956_(_05565_, _05564_, _02089_);
    or _11957_(_00083_, _05565_, _05550_);
    and _11958_(_05566_, _02090_, base[12]);
    nor _11959_(_05567_, _02095_, _01934_);
    or _11960_(_05568_, _01954_, modulus[11]);
    or _11961_(_05569_, _05553_, _01956_);
    and _11962_(_05570_, _05569_, _05568_);
    or _11963_(_05571_, _05537_, _01966_);
    and _11964_(_05572_, _05571_, _05570_);
    or _11965_(_05574_, _05506_, _01991_);
    and _11966_(_05575_, _05574_, _05572_);
    xnor _11967_(_05576_, _05575_, _01943_);
    nor _11968_(_05577_, _05576_, _02079_);
    or _11969_(_05578_, _05577_, _05567_);
    and _11970_(_05579_, _05578_, _02084_);
    and _11971_(_05580_, _05579_, rsa_active);
    and _11972_(_05581_, _05580_, _02093_);
    and _11973_(_05582_, _01160_, message[12]);
    or _11974_(_05583_, _05582_, _05581_);
    and _11975_(_05585_, _05583_, _02089_);
    or _11976_(_00084_, _05585_, _05566_);
    and _11977_(_05586_, _02090_, base[13]);
    nor _11978_(_05587_, _02095_, _01927_);
    or _11979_(_05588_, _01934_, modulus[12]);
    or _11980_(_05589_, _05575_, _01943_);
    and _11981_(_05590_, _05589_, _05588_);
    xnor _11982_(_05591_, _05590_, _01930_);
    nor _11983_(_05592_, _05591_, _02079_);
    or _11984_(_05593_, _05592_, _05587_);
    and _11985_(_05595_, _05593_, _02084_);
    and _11986_(_05596_, _05595_, rsa_active);
    and _11987_(_05597_, _05596_, _02093_);
    and _11988_(_05598_, _01160_, message[13]);
    or _11989_(_05599_, _05598_, _05597_);
    and _11990_(_05600_, _05599_, _02089_);
    or _11991_(_00085_, _05600_, _05586_);
    and _11992_(_05601_, _02090_, base[14]);
    nor _11993_(_05602_, _02095_, _01915_);
    or _11994_(_05603_, _01927_, modulus[13]);
    or _11995_(_05605_, _05588_, _01930_);
    and _11996_(_05606_, _05605_, _05603_);
    not _11997_(_05607_, _01944_);
    or _11998_(_05608_, _05575_, _05607_);
    and _11999_(_05609_, _05608_, _05606_);
    xnor _12000_(_05610_, _05609_, _01920_);
    nor _12001_(_05611_, _05610_, _02079_);
    or _12002_(_05612_, _05611_, _05602_);
    and _12003_(_05613_, _05612_, _02084_);
    and _12004_(_05614_, _05613_, rsa_active);
    and _12005_(_05616_, _05614_, _02093_);
    and _12006_(_05617_, _01160_, message[14]);
    or _12007_(_05618_, _05617_, _05616_);
    and _12008_(_05619_, _05618_, _02089_);
    or _12009_(_00086_, _05619_, _05601_);
    and _12010_(_05620_, _02090_, base[15]);
    nor _12011_(_05621_, _02095_, _01910_);
    or _12012_(_05622_, _01915_, modulus[14]);
    or _12013_(_05623_, _05609_, _01920_);
    and _12014_(_05624_, _05623_, _05622_);
    xor _12015_(_05626_, _05624_, _01911_);
    and _12016_(_05627_, _05626_, _02095_);
    or _12017_(_05628_, _05627_, _05621_);
    and _12018_(_05629_, _05628_, _02084_);
    and _12019_(_05630_, _05629_, rsa_active);
    and _12020_(_05631_, _05630_, _02093_);
    and _12021_(_05632_, _01160_, message[15]);
    or _12022_(_05633_, _05632_, _05631_);
    and _12023_(_05634_, _05633_, _02089_);
    or _12024_(_00087_, _05634_, _05620_);
    and _12025_(_05636_, _02090_, exp_counter[0]);
    and _12026_(_05637_, _02084_, exp_counter[1]);
    and _12027_(_05638_, _05637_, rsa_active);
    and _12028_(_05639_, _05638_, _02093_);
    and _12029_(_05640_, _01160_, exponent[0]);
    or _12030_(_05641_, _05640_, _05639_);
    and _12031_(_05642_, _05641_, _02089_);
    or _12032_(_00088_, _05642_, _05636_);
    and _12033_(_05643_, _02090_, exp_counter[1]);
    and _12034_(_05644_, _02084_, exp_counter[2]);
    and _12035_(_05646_, _05644_, rsa_active);
    and _12036_(_05647_, _05646_, _02093_);
    and _12037_(_05648_, _01160_, exponent[1]);
    or _12038_(_05649_, _05648_, _05647_);
    and _12039_(_05650_, _05649_, _02089_);
    or _12040_(_00089_, _05650_, _05643_);
    and _12041_(_05651_, _02090_, exp_counter[2]);
    and _12042_(_05652_, _02084_, exp_counter[3]);
    and _12043_(_05653_, _05652_, rsa_active);
    and _12044_(_05654_, _05653_, _02093_);
    and _12045_(_05656_, _01160_, exponent[2]);
    or _12046_(_05657_, _05656_, _05654_);
    and _12047_(_05658_, _05657_, _02089_);
    or _12048_(_00090_, _05658_, _05651_);
    and _12049_(_05659_, _02090_, exp_counter[3]);
    and _12050_(_05660_, _01160_, exponent[3]);
    and _12051_(_05661_, _05660_, _02089_);
    or _12052_(_00091_, _05661_, _05659_);
    and _12053_(_05662_, _02108_, result[0]);
    and _12054_(_05663_, _02107_, accumulator[0]);
    or _12055_(_00092_, _05663_, _05662_);
    and _12056_(_05665_, _02108_, result[1]);
    and _12057_(_05666_, _02107_, accumulator[1]);
    or _12058_(_00093_, _05666_, _05665_);
    and _12059_(_05667_, _02108_, result[2]);
    and _12060_(_05668_, _02107_, accumulator[2]);
    or _12061_(_00094_, _05668_, _05667_);
    and _12062_(_05669_, _02108_, result[3]);
    and _12063_(_05670_, _02107_, accumulator[3]);
    or _12064_(_00095_, _05670_, _05669_);
    and _12065_(_05672_, _02108_, result[4]);
    and _12066_(_05673_, _02107_, accumulator[4]);
    or _12067_(_00096_, _05673_, _05672_);
    and _12068_(_05674_, _02108_, result[5]);
    and _12069_(_05675_, _02107_, accumulator[5]);
    or _12070_(_00097_, _05675_, _05674_);
    and _12071_(_05676_, _02108_, result[6]);
    and _12072_(_05677_, _02107_, accumulator[6]);
    or _12073_(_00098_, _05677_, _05676_);
    and _12074_(_05678_, _02108_, result[7]);
    and _12075_(_05680_, _02107_, accumulator[7]);
    or _12076_(_00099_, _05680_, _05678_);
    and _12077_(_05681_, _02108_, result[8]);
    and _12078_(_05682_, _02107_, accumulator[8]);
    or _12079_(_00100_, _05682_, _05681_);
    and _12080_(_05683_, _02108_, result[9]);
    and _12081_(_05684_, _02107_, accumulator[9]);
    or _12082_(_00101_, _05684_, _05683_);
    and _12083_(_05685_, _02108_, result[10]);
    and _12084_(_05686_, _02107_, accumulator[10]);
    or _12085_(_00102_, _05686_, _05685_);
    and _12086_(_05688_, _02108_, result[11]);
    and _12087_(_05689_, _02107_, accumulator[11]);
    or _12088_(_00103_, _05689_, _05688_);
    and _12089_(_05690_, _02108_, result[12]);
    and _12090_(_05691_, _02107_, accumulator[12]);
    or _12091_(_00104_, _05691_, _05690_);
    and _12092_(_05692_, _02108_, result[13]);
    and _12093_(_05693_, _02107_, accumulator[13]);
    or _12094_(_00105_, _05693_, _05692_);
    and _12095_(_05695_, _02108_, result[14]);
    and _12096_(_05696_, _02107_, accumulator[14]);
    or _12097_(_00106_, _05696_, _05695_);
    and _12098_(_05697_, _02108_, result[15]);
    and _12099_(_05698_, _02107_, accumulator[15]);
    or _12100_(_00107_, _05698_, _05697_);
    nor _12101_(_05699_, _02082_, _01149_);
    or _12102_(_00000_, _05699_, _01160_);
    not _12103_(_00002_, rst);
    not _12104_(_00003_, rst);
    not _12105_(_00004_, rst);
    not _12106_(_00005_, rst);
    not _12107_(_00006_, rst);
    not _12108_(_00007_, rst);
    not _12109_(_00008_, rst);
    not _12110_(_00009_, rst);
    not _12111_(_00010_, rst);
    not _12112_(_00011_, rst);
    not _12113_(_00012_, rst);
    not _12114_(_00013_, rst);
    not _12115_(_00014_, rst);
    not _12116_(_00015_, rst);
    not _12117_(_00016_, rst);
    not _12118_(_00017_, rst);
    not _12119_(_00018_, rst);
    not _12120_(_00019_, rst);
    not _12121_(_00020_, rst);
    not _12122_(_00021_, rst);
    not _12123_(_00022_, rst);
    not _12124_(_00023_, rst);
    not _12125_(_00024_, rst);
    not _12126_(_00025_, rst);
    not _12127_(_00026_, rst);
    not _12128_(_00027_, rst);
    not _12129_(_00028_, rst);
    not _12130_(_00029_, rst);
    not _12131_(_00030_, rst);
    not _12132_(_00031_, rst);
    not _12133_(_00032_, rst);
    not _12134_(_00033_, rst);
    not _12135_(_00034_, rst);
    not _12136_(_00035_, rst);
    not _12137_(_00036_, rst);
    not _12138_(_00037_, rst);
    not _12139_(_00038_, rst);
    not _12140_(_00039_, rst);
    not _12141_(_00040_, rst);
    not _12142_(_00041_, rst);
    not _12143_(_00042_, rst);
    not _12144_(_00043_, rst);
    not _12145_(_00044_, rst);
    not _12146_(_00045_, rst);
    not _12147_(_00046_, rst);
    not _12148_(_00047_, rst);
    not _12149_(_00048_, rst);
    not _12150_(_00049_, rst);
    not _12151_(_00050_, rst);
    not _12152_(_00051_, rst);
    not _12153_(_00052_, rst);
    not _12154_(_00053_, rst);
    not _12155_(_00054_, rst);
    dff _12156_(.RN(_00001_), .SN(1'b1), .CK(clk), .D(_00055_), .Q(base[0]));
    dff _12157_(.RN(_00002_), .SN(1'b1), .CK(clk), .D(_00056_), .Q(rsa_done));
    dff _12158_(.RN(_00003_), .SN(1'b1), .CK(clk), .D(_00057_), .Q(accumulator[0]));
    dff _12159_(.RN(_00004_), .SN(1'b1), .CK(clk), .D(_00058_), .Q(accumulator[1]));
    dff _12160_(.RN(_00005_), .SN(1'b1), .CK(clk), .D(_00059_), .Q(accumulator[2]));
    dff _12161_(.RN(_00006_), .SN(1'b1), .CK(clk), .D(_00060_), .Q(accumulator[3]));
    dff _12162_(.RN(_00007_), .SN(1'b1), .CK(clk), .D(_00061_), .Q(accumulator[4]));
    dff _12163_(.RN(_00008_), .SN(1'b1), .CK(clk), .D(_00062_), .Q(accumulator[5]));
    dff _12164_(.RN(_00009_), .SN(1'b1), .CK(clk), .D(_00063_), .Q(accumulator[6]));
    dff _12165_(.RN(_00010_), .SN(1'b1), .CK(clk), .D(_00064_), .Q(accumulator[7]));
    dff _12166_(.RN(_00011_), .SN(1'b1), .CK(clk), .D(_00065_), .Q(accumulator[8]));
    dff _12167_(.RN(_00012_), .SN(1'b1), .CK(clk), .D(_00066_), .Q(accumulator[9]));
    dff _12168_(.RN(_00013_), .SN(1'b1), .CK(clk), .D(_00067_), .Q(accumulator[10]));
    dff _12169_(.RN(_00014_), .SN(1'b1), .CK(clk), .D(_00068_), .Q(accumulator[11]));
    dff _12170_(.RN(_00015_), .SN(1'b1), .CK(clk), .D(_00069_), .Q(accumulator[12]));
    dff _12171_(.RN(_00016_), .SN(1'b1), .CK(clk), .D(_00070_), .Q(accumulator[13]));
    dff _12172_(.RN(_00017_), .SN(1'b1), .CK(clk), .D(_00071_), .Q(accumulator[14]));
    dff _12173_(.RN(_00018_), .SN(1'b1), .CK(clk), .D(_00072_), .Q(accumulator[15]));
    dff _12174_(.RN(_00019_), .SN(1'b1), .CK(clk), .D(_00073_), .Q(base[1]));
    dff _12175_(.RN(_00020_), .SN(1'b1), .CK(clk), .D(_00074_), .Q(base[2]));
    dff _12176_(.RN(_00021_), .SN(1'b1), .CK(clk), .D(_00075_), .Q(base[3]));
    dff _12177_(.RN(_00022_), .SN(1'b1), .CK(clk), .D(_00076_), .Q(base[4]));
    dff _12178_(.RN(_00023_), .SN(1'b1), .CK(clk), .D(_00077_), .Q(base[5]));
    dff _12179_(.RN(_00024_), .SN(1'b1), .CK(clk), .D(_00078_), .Q(base[6]));
    dff _12180_(.RN(_00025_), .SN(1'b1), .CK(clk), .D(_00079_), .Q(base[7]));
    dff _12181_(.RN(_00026_), .SN(1'b1), .CK(clk), .D(_00080_), .Q(base[8]));
    dff _12182_(.RN(_00027_), .SN(1'b1), .CK(clk), .D(_00081_), .Q(base[9]));
    dff _12183_(.RN(_00028_), .SN(1'b1), .CK(clk), .D(_00082_), .Q(base[10]));
    dff _12184_(.RN(_00029_), .SN(1'b1), .CK(clk), .D(_00083_), .Q(base[11]));
    dff _12185_(.RN(_00030_), .SN(1'b1), .CK(clk), .D(_00084_), .Q(base[12]));
    dff _12186_(.RN(_00031_), .SN(1'b1), .CK(clk), .D(_00085_), .Q(base[13]));
    dff _12187_(.RN(_00032_), .SN(1'b1), .CK(clk), .D(_00086_), .Q(base[14]));
    dff _12188_(.RN(_00033_), .SN(1'b1), .CK(clk), .D(_00087_), .Q(base[15]));
    dff _12189_(.RN(_00034_), .SN(1'b1), .CK(clk), .D(_00088_), .Q(exp_counter[0]));
    dff _12190_(.RN(_00035_), .SN(1'b1), .CK(clk), .D(_00089_), .Q(exp_counter[1]));
    dff _12191_(.RN(_00036_), .SN(1'b1), .CK(clk), .D(_00090_), .Q(exp_counter[2]));
    dff _12192_(.RN(_00037_), .SN(1'b1), .CK(clk), .D(_00091_), .Q(exp_counter[3]));
    dff _12193_(.RN(_00038_), .SN(1'b1), .CK(clk), .D(_00000_), .Q(rsa_active));
    dff _12194_(.RN(_00039_), .SN(1'b1), .CK(clk), .D(_00092_), .Q(result[0]));
    dff _12195_(.RN(_00040_), .SN(1'b1), .CK(clk), .D(_00093_), .Q(result[1]));
    dff _12196_(.RN(_00041_), .SN(1'b1), .CK(clk), .D(_00094_), .Q(result[2]));
    dff _12197_(.RN(_00042_), .SN(1'b1), .CK(clk), .D(_00095_), .Q(result[3]));
    dff _12198_(.RN(_00043_), .SN(1'b1), .CK(clk), .D(_00096_), .Q(result[4]));
    dff _12199_(.RN(_00044_), .SN(1'b1), .CK(clk), .D(_00097_), .Q(result[5]));
    dff _12200_(.RN(_00045_), .SN(1'b1), .CK(clk), .D(_00098_), .Q(result[6]));
    dff _12201_(.RN(_00046_), .SN(1'b1), .CK(clk), .D(_00099_), .Q(result[7]));
    dff _12202_(.RN(_00047_), .SN(1'b1), .CK(clk), .D(_00100_), .Q(result[8]));
    dff _12203_(.RN(_00048_), .SN(1'b1), .CK(clk), .D(_00101_), .Q(result[9]));
    dff _12204_(.RN(_00049_), .SN(1'b1), .CK(clk), .D(_00102_), .Q(result[10]));
    dff _12205_(.RN(_00050_), .SN(1'b1), .CK(clk), .D(_00103_), .Q(result[11]));
    dff _12206_(.RN(_00051_), .SN(1'b1), .CK(clk), .D(_00104_), .Q(result[12]));
    dff _12207_(.RN(_00052_), .SN(1'b1), .CK(clk), .D(_00105_), .Q(result[13]));
    dff _12208_(.RN(_00053_), .SN(1'b1), .CK(clk), .D(_00106_), .Q(result[14]));
    dff _12209_(.RN(_00054_), .SN(1'b1), .CK(clk), .D(_00107_), .Q(result[15]));
endmodule