module trojan0_crypto0_host_0000(clk, rst, plaintext, cipher_key, encrypt_start, ciphertext, encrypt_done);
  wire _0000_;
  wire _0001_;
  wire _0002_;
  wire _0003_;
  wire _0004_;
  wire _0005_;
  wire _0006_;
  wire _0007_;
  wire _0008_;
  wire _0009_;
  wire _0010_;
  wire _0011_;
  wire _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  wire _0514_;
  wire _0515_;
  wire _0516_;
  wire _0517_;
  wire _0518_;
  wire _0519_;
  wire _0520_;
  wire _0521_;
  wire _0522_;
  wire _0523_;
  wire _0524_;
  wire _0525_;
  wire _0526_;
  wire _0527_;
  wire _0528_;
  wire _0529_;
  wire _0530_;
  wire _0531_;
  wire _0532_;
  wire _0533_;
  wire _0534_;
  wire _0535_;
  wire _0536_;
  wire _0537_;
  wire _0538_;
  wire _0539_;
  wire _0540_;
  wire _0541_;
  wire _0542_;
  wire _0543_;
  wire _0544_;
  wire _0545_;
  wire _0546_;
  wire _0547_;
  wire _0548_;
  wire _0549_;
  wire _0550_;
  wire _0551_;
  wire _0552_;
  wire _0553_;
  wire _0554_;
  wire _0555_;
  wire _0556_;
  wire _0557_;
  wire _0558_;
  wire _0559_;
  wire _0560_;
  wire _0561_;
  wire _0562_;
  wire _0563_;
  wire _0564_;
  wire _0565_;
  wire _0566_;
  wire _0567_;
  wire _0568_;
  wire _0569_;
  wire _0570_;
  wire _0571_;
  wire _0572_;
  wire _0573_;
  wire _0574_;
  wire _0575_;
  wire _0576_;
  wire _0577_;
  wire _0578_;
  wire _0579_;
  wire _0580_;
  wire _0581_;
  wire _0582_;
  wire _0583_;
  wire _0584_;
  wire _0585_;
  wire _0586_;
  wire _0587_;
  wire _0588_;
  wire _0589_;
  wire _0590_;
  wire _0591_;
  wire _0592_;
  wire _0593_;
  wire _0594_;
  wire _0595_;
  wire _0596_;
  wire _0597_;
  wire _0598_;
  wire _0599_;
  wire _0600_;
  wire _0601_;
  wire _0602_;
  wire _0603_;
  wire _0604_;
  wire _0605_;
  wire _0606_;
  wire _0607_;
  wire _0608_;
  wire _0609_;
  wire _0610_;
  wire _0611_;
  wire _0612_;
  wire _0613_;
  wire _0614_;
  wire _0615_;
  wire _0616_;
  wire _0617_;
  wire _0618_;
  wire _0619_;
  wire _0620_;
  wire _0621_;
  wire _0622_;
  wire _0623_;
  wire _0624_;
  wire _0625_;
  wire _0626_;
  wire _0627_;
  wire _0628_;
  wire _0629_;
  wire _0630_;
  wire _0631_;
  wire _0632_;
  wire _0633_;
  wire _0634_;
  wire _0635_;
  wire _0636_;
  wire _0637_;
  wire _0638_;
  wire _0639_;
  wire _0640_;
  wire _0641_;
  wire _0642_;
  wire _0643_;
  wire _0644_;
  wire _0645_;
  wire _0646_;
  wire _0647_;
  wire _0648_;
  wire _0649_;
  wire _0650_;
  wire _0651_;
  wire _0652_;
  wire _0653_;
  wire _0654_;
  wire _0655_;
  wire _0656_;
  wire _0657_;
  wire _0658_;
  wire _0659_;
  wire _0660_;
  wire _0661_;
  wire _0662_;
  wire _0663_;
  wire _0664_;
  wire _0665_;
  wire _0666_;
  wire _0667_;
  wire _0668_;
  wire _0669_;
  wire _0670_;
  wire _0671_;
  wire _0672_;
  wire _0673_;
  wire _0674_;
  wire _0675_;
  wire _0676_;
  wire _0677_;
  wire _0678_;
  wire _0679_;
  wire _0680_;
  wire _0681_;
  wire _0682_;
  wire _0683_;
  wire _0684_;
  wire _0685_;
  wire _0686_;
  wire _0687_;
  wire _0688_;
  wire _0689_;
  wire _0690_;
  wire _0691_;
  wire _0692_;
  wire _0693_;
  wire _0694_;
  wire _0695_;
  wire _0696_;
  wire _0697_;
  wire _0698_;
  wire _0699_;
  wire _0700_;
  wire _0701_;
  wire _0702_;
  wire _0703_;
  wire _0704_;
  wire _0705_;
  wire _0706_;
  wire _0707_;
  wire _0708_;
  wire _0709_;
  wire _0710_;
  wire _0711_;
  wire _0712_;
  wire _0713_;
  wire _0714_;
  wire _0715_;
  wire _0716_;
  wire _0717_;
  wire _0718_;
  wire _0719_;
  wire _0720_;
  wire _0721_;
  wire _0722_;
  wire _0723_;
  wire _0724_;
  wire _0725_;
  wire _0726_;
  wire _0727_;
  wire _0728_;
  wire _0729_;
  wire _0730_;
  wire _0731_;
  wire _0732_;
  wire _0733_;
  wire _0734_;
  wire _0735_;
  wire _0736_;
  wire _0737_;
  wire _0738_;
  wire _0739_;
  wire _0740_;
  wire _0741_;
  wire _0742_;
  wire _0743_;
  wire _0744_;
  wire _0745_;
  wire _0746_;
  wire _0747_;
  wire _0748_;
  wire _0749_;
  wire _0750_;
  wire _0751_;
  wire _0752_;
  wire _0753_;
  wire _0754_;
  wire _0755_;
  wire _0756_;
  wire _0757_;
  wire _0758_;
  wire _0759_;
  wire _0760_;
  wire _0761_;
  wire _0762_;
  wire _0763_;
  wire _0764_;
  wire _0765_;
  wire _0766_;
  wire _0767_;
  wire _0768_;
  wire _0769_;
  wire _0770_;
  wire _0771_;
  wire _0772_;
  wire _0773_;
  wire _0774_;
  wire _0775_;
  wire _0776_;
  wire _0777_;
  wire _0778_;
  wire _0779_;
  wire _0780_;
  wire _0781_;
  wire _0782_;
  wire _0783_;
  wire _0784_;
  wire _0785_;
  wire _0786_;
  wire _0787_;
  wire _0788_;
  wire _0789_;
  wire _0790_;
  wire _0791_;
  wire _0792_;
  wire _0793_;
  wire _0794_;
  wire _0795_;
  wire _0796_;
  wire _0797_;
  wire _0798_;
  wire _0799_;
  wire _0800_;
  wire _0801_;
  wire _0802_;
  wire _0803_;
  wire _0804_;
  wire _0805_;
  wire _0806_;
  wire _0807_;
  wire _0808_;
  wire _0809_;
  wire _0810_;
  wire _0811_;
  wire _0812_;
  wire _0813_;
  wire _0814_;
  wire _0815_;
  wire _0816_;
  wire _0817_;
  wire _0818_;
  wire _0819_;
  wire _0820_;
  wire _0821_;
  wire _0822_;
  wire _0823_;
  wire _0824_;
  wire _0825_;
  wire _0826_;
  wire _0827_;
  wire _0828_;
  wire _0829_;
  wire _0830_;
  wire _0831_;
  wire _0832_;
  wire _0833_;
  wire _0834_;
  wire _0835_;
  wire _0836_;
  wire _0837_;
  wire _0838_;
  wire _0839_;
  wire _0840_;
  wire _0841_;
  wire _0842_;
  wire _0843_;
  wire _0844_;
  wire _0845_;
  wire _0846_;
  wire _0847_;
  wire _0848_;
  wire _0849_;
  wire _0850_;
  wire _0851_;
  wire _0852_;
  wire _0853_;
  wire _0854_;
  wire _0855_;
  wire _0856_;
  wire _0857_;
  wire _0858_;
  wire _0859_;
  wire _0860_;
  wire _0861_;
  wire _0862_;
  wire _0863_;
  wire _0864_;
  wire _0865_;
  wire _0866_;
  wire _0867_;
  wire _0868_;
  wire _0869_;
  wire _0870_;
  wire _0871_;
  wire _0872_;
  wire _0873_;
  wire _0874_;
  wire _0875_;
  wire _0876_;
  wire _0877_;
  wire _0878_;
  wire _0879_;
  wire _0880_;
  wire _0881_;
  wire _0882_;
  wire _0883_;
  wire _0884_;
  wire _0885_;
  wire _0886_;
  wire _0887_;
  wire _0888_;
  wire _0889_;
  wire _0890_;
  wire _0891_;
  wire _0892_;
  wire _0893_;
  wire _0894_;
  wire _0895_;
  wire _0896_;
  wire _0897_;
  wire _0898_;
  wire _0899_;
  wire _0900_;
  wire _0901_;
  wire _0902_;
  wire _0903_;
  wire _0904_;
  wire _0905_;
  wire _0906_;
  wire _0907_;
  wire _0908_;
  wire _0909_;
  wire _0910_;
  wire _0911_;
  wire _0912_;
  wire _0913_;
  wire _0914_;
  wire _0915_;
  wire _0916_;
  wire _0917_;
  wire _0918_;
  wire _0919_;
  wire _0920_;
  wire _0921_;
  wire _0922_;
  wire _0923_;
  wire _0924_;
  wire _0925_;
  wire _0926_;
  wire _0927_;
  wire _0928_;
  wire _0929_;
  wire _0930_;
  wire _0931_;
  wire _0932_;
  wire _0933_;
  wire _0934_;
  wire _0935_;
  wire _0936_;
  wire _0937_;
  wire _0938_;
  wire _0939_;
  wire _0940_;
  wire _0941_;
  wire _0942_;
  wire _0943_;
  wire _0944_;
  wire _0945_;
  wire _0946_;
  wire _0947_;
  wire _0948_;
  wire _0949_;
  wire _0950_;
  wire _0951_;
  wire _0952_;
  wire _0953_;
  wire _0954_;
  wire _0955_;
  wire _0956_;
  wire _0957_;
  wire _0958_;
  wire _0959_;
  wire _0960_;
  wire _0961_;
  wire _0962_;
  wire _0963_;
  wire _0964_;
  wire _0965_;
  wire _0966_;
  wire _0967_;
  wire _0968_;
  wire _0969_;
  wire _0970_;
  wire _0971_;
  wire _0972_;
  wire _0973_;
  wire _0974_;
  wire _0975_;
  wire _0976_;
  wire _0977_;
  wire _0978_;
  wire _0979_;
  wire _0980_;
  wire _0981_;
  wire _0982_;
  wire _0983_;
  wire _0984_;
  wire _0985_;
  wire _0986_;
  wire _0987_;
  wire _0988_;
  wire _0989_;
  wire _0990_;
  wire _0991_;
  wire _0992_;
  wire _0993_;
  wire _0994_;
  wire _0995_;
  wire _0996_;
  wire _0997_;
  wire _0998_;
  wire _0999_;
  wire _1000_;
  wire _1001_;
  wire _1002_;
  wire _1003_;
  wire _1004_;
  wire _1005_;
  wire _1006_;
  wire _1007_;
  wire _1008_;
  wire _1009_;
  wire _1010_;
  wire _1011_;
  wire _1012_;
  wire _1013_;
  wire _1014_;
  wire _1015_;
  wire _1016_;
  wire _1017_;
  wire _1018_;
  wire _1019_;
  wire _1020_;
  wire _1021_;
  wire _1022_;
  wire _1023_;
  wire _1024_;
  wire _1025_;
  wire _1026_;
  wire _1027_;
  wire _1028_;
  wire _1029_;
  wire _1030_;
  wire _1031_;
  wire _1032_;
  wire _1033_;
  wire _1034_;
  wire _1035_;
  wire _1036_;
  wire _1037_;
  wire _1038_;
  wire _1039_;
  wire _1040_;
  wire _1041_;
  wire _1042_;
  wire _1043_;
  wire _1044_;
  wire _1045_;
  wire _1046_;
  wire _1047_;
  wire _1048_;
  wire _1049_;
  wire _1050_;
  wire _1051_;
  wire _1052_;
  wire _1053_;
  wire _1054_;
  wire _1055_;
  wire _1056_;
  wire _1057_;
  wire _1058_;
  wire _1059_;
  wire _1060_;
  wire _1061_;
  wire _1062_;
  wire _1063_;
  wire _1064_;
  wire _1065_;
  wire _1066_;
  wire _1067_;
  wire _1068_;
  wire _1069_;
  wire _1070_;
  wire _1071_;
  wire _1072_;
  wire _1073_;
  wire _1074_;
  wire _1075_;
  wire _1076_;
  wire _1077_;
  wire _1078_;
  wire _1079_;
  wire _1080_;
  wire _1081_;
  wire _1082_;
  wire _1083_;
  wire _1084_;
  wire _1085_;
  wire _1086_;
  wire _1087_;
  wire _1088_;
  wire _1089_;
  wire _1090_;
  wire _1091_;
  wire _1092_;
  wire _1093_;
  wire _1094_;
  wire _1095_;
  wire _1096_;
  wire _1097_;
  wire _1098_;
  wire _1099_;
  wire _1100_;
  wire _1101_;
  wire _1102_;
  wire _1103_;
  wire _1104_;
  wire _1105_;
  wire _1106_;
  wire _1107_;
  wire _1108_;
  wire _1109_;
  wire _1110_;
  wire _1111_;
  wire _1112_;
  wire _1113_;
  wire _1114_;
  wire _1115_;
  wire _1116_;
  wire _1117_;
  wire _1118_;
  wire _1119_;
  wire _1120_;
  wire _1121_;
  wire _1122_;
  wire _1123_;
  wire _1124_;
  wire _1125_;
  wire _1126_;
  wire _1127_;
  wire _1128_;
  wire _1129_;
  wire _1130_;
  wire _1131_;
  wire _1132_;
  wire _1133_;
  wire _1134_;
  wire _1135_;
  wire _1136_;
  wire _1137_;
  wire _1138_;
  wire _1139_;
  wire _1140_;
  wire _1141_;
  wire _1142_;
  wire _1143_;
  wire _1144_;
  wire _1145_;
  wire _1146_;
  wire _1147_;
  wire _1148_;
  wire _1149_;
  wire _1150_;
  wire _1151_;
  wire _1152_;
  wire _1153_;
  wire _1154_;
  wire _1155_;
  wire _1156_;
  wire _1157_;
  wire _1158_;
  wire _1159_;
  wire _1160_;
  wire _1161_;
  wire _1162_;
  wire _1163_;
  wire _1164_;
  wire _1165_;
  wire _1166_;
  wire _1167_;
  wire _1168_;
  wire _1169_;
  wire _1170_;
  wire _1171_;
  wire _1172_;
  wire _1173_;
  wire _1174_;
  wire _1175_;
  wire _1176_;
  wire _1177_;
  wire _1178_;
  wire _1179_;
  wire _1180_;
  wire _1181_;
  wire _1182_;
  wire _1183_;
  wire _1184_;
  wire _1185_;
  wire _1186_;
  wire _1187_;
  wire _1188_;
  wire _1189_;
  wire _1190_;
  wire _1191_;
  wire _1192_;
  wire _1193_;
  wire _1194_;
  wire _1195_;
  wire _1196_;
  wire _1197_;
  wire _1198_;
  wire _1199_;
  wire _1200_;
  wire _1201_;
  wire _1202_;
  wire _1203_;
  wire _1204_;
  wire _1205_;
  wire _1206_;
  wire _1207_;
  wire _1208_;
  wire _1209_;
  wire _1210_;
  wire _1211_;
  wire _1212_;
  wire _1213_;
  wire _1214_;
  wire _1215_;
  wire _1216_;
  wire _1217_;
  wire _1218_;
  wire _1219_;
  wire _1220_;
  wire _1221_;
  wire _1222_;
  wire _1223_;
  wire _1224_;
  wire _1225_;
  wire _1226_;
  wire _1227_;
  wire _1228_;
  wire _1229_;
  wire _1230_;
  wire _1231_;
  wire _1232_;
  wire _1233_;
  wire _1234_;
  wire _1235_;
  wire _1236_;
  wire _1237_;
  wire _1238_;
  wire _1239_;
  wire _1240_;
  wire _1241_;
  wire _1242_;
  wire _1243_;
  wire _1244_;
  wire _1245_;
  wire _1246_;
  wire _1247_;
  wire _1248_;
  wire _1249_;
  wire _1250_;
  wire _1251_;
  wire _1252_;
  wire _1253_;
  wire _1254_;
  wire _1255_;
  wire _1256_;
  wire _1257_;
  wire _1258_;
  wire _1259_;
  wire _1260_;
  wire _1261_;
  wire _1262_;
  wire _1263_;
  wire _1264_;
  wire _1265_;
  wire _1266_;
  wire _1267_;
  wire _1268_;
  wire _1269_;
  wire _1270_;
  wire _1271_;
  wire _1272_;
  wire _1273_;
  wire _1274_;
  wire _1275_;
  wire _1276_;
  wire _1277_;
  wire _1278_;
  wire _1279_;
  wire _1280_;
  wire _1281_;
  wire _1282_;
  wire _1283_;
  wire _1284_;
  wire _1285_;
  wire _1286_;
  wire _1287_;
  wire _1288_;
  wire _1289_;
  wire _1290_;
  wire _1291_;
  wire _1292_;
  wire _1293_;
  wire _1294_;
  wire _1295_;
  wire _1296_;
  wire _1297_;
  wire _1298_;
  wire _1299_;
  wire _1300_;
  wire _1301_;
  wire _1302_;
  wire _1303_;
  wire _1304_;
  wire _1305_;
  wire _1306_;
  wire _1307_;
  wire _1308_;
  wire _1309_;
  wire _1310_;
  wire _1311_;
  wire _1312_;
  wire _1313_;
  wire _1314_;
  wire _1315_;
  wire _1316_;
  wire _1317_;
  wire _1318_;
  wire _1319_;
  wire _1320_;
  wire _1321_;
  wire _1322_;
  wire _1323_;
  wire _1324_;
  wire _1325_;
  wire _1326_;
  wire _1327_;
  wire _1328_;
  wire _1329_;
  wire _1330_;
  wire _1331_;
  wire _1332_;
  wire _1333_;
  wire _1334_;
  wire _1335_;
  wire _1336_;
  wire _1337_;
  wire _1338_;
  wire _1339_;
  wire _1340_;
  wire _1341_;
  wire _1342_;
  wire _1343_;
  wire _1344_;
  wire _1345_;
  wire _1346_;
  wire _1347_;
  wire _1348_;
  wire _1349_;
  wire _1350_;
  wire _1351_;
  wire _1352_;
  wire _1353_;
  wire _1354_;
  wire _1355_;
  wire _1356_;
  wire _1357_;
  wire _1358_;
  wire _1359_;
  wire _1360_;
  wire _1361_;
  wire _1362_;
  wire _1363_;
  wire _1364_;
  wire _1365_;
  wire _1366_;
  wire _1367_;
  wire _1368_;
  wire _1369_;
  wire _1370_;
  wire _1371_;
  wire _1372_;
  wire _1373_;
  wire _1374_;
  wire _1375_;
  wire _1376_;
  wire _1377_;
  wire _1378_;
  wire _1379_;
  wire _1380_;
  wire _1381_;
  wire _1382_;
  wire _1383_;
  wire _1384_;
  wire _1385_;
  wire _1386_;
  wire _1387_;
  wire _1388_;
  wire _1389_;
  wire _1390_;
  wire _1391_;
  wire _1392_;
  wire _1393_;
  wire _1394_;
  wire _1395_;
  wire _1396_;
  wire _1397_;
  wire _1398_;
  wire _1399_;
  wire _1400_;
  wire _1401_;
  wire _1402_;
  wire _1403_;
  wire _1404_;
  wire _1405_;
  wire _1406_;
  wire _1407_;
  wire _1408_;
  wire _1409_;
  wire _1410_;
  wire _1411_;
  wire _1412_;
  wire _1413_;
  wire _1414_;
  wire _1415_;
  wire _1416_;
  wire _1417_;
  wire _1418_;
  wire _1419_;
  wire _1420_;
  wire _1421_;
  wire _1422_;
  wire _1423_;
  wire _1424_;
  wire _1425_;
  wire _1426_;
  wire _1427_;
  wire _1428_;
  wire _1429_;
  wire _1430_;
  wire _1431_;
  wire _1432_;
  wire _1433_;
  wire _1434_;
  wire _1435_;
  wire _1436_;
  wire _1437_;
  wire _1438_;
  wire _1439_;
  wire _1440_;
  wire _1441_;
  wire _1442_;
  wire _1443_;
  wire _1444_;
  wire _1445_;
  wire _1446_;
  wire _1447_;
  wire _1448_;
  wire _1449_;
  wire _1450_;
  wire _1451_;
  wire _1452_;
  wire _1453_;
  wire _1454_;
  wire _1455_;
  wire _1456_;
  wire _1457_;
  wire _1458_;
  wire _1459_;
  wire _1460_;
  wire _1461_;
  wire _1462_;
  wire _1463_;
  wire _1464_;
  wire _1465_;
  wire _1466_;
  wire _1467_;
  wire _1468_;
  wire _1469_;
  wire _1470_;
  wire _1471_;
  wire _1472_;
  wire _1473_;
  wire _1474_;
  wire _1475_;
  wire _1476_;
  wire _1477_;
  wire _1478_;
  wire _1479_;
  wire _1480_;
  wire _1481_;
  wire _1482_;
  wire _1483_;
  wire _1484_;
  wire _1485_;
  wire _1486_;
  wire _1487_;
  wire _1488_;
  wire _1489_;
  wire _1490_;
  wire _1491_;
  wire _1492_;
  wire _1493_;
  wire _1494_;
  wire _1495_;
  wire _1496_;
  wire _1497_;
  wire _1498_;
  wire _1499_;
  wire _1500_;
  wire _1501_;
  wire _1502_;
  wire _1503_;
  wire _1504_;
  wire _1505_;
  wire _1506_;
  wire _1507_;
  wire _1508_;
  wire _1509_;
  wire _1510_;
  wire _1511_;
  wire _1512_;
  wire _1513_;
  wire _1514_;
  wire _1515_;
  wire _1516_;
  wire _1517_;
  wire _1518_;
  wire _1519_;
  wire _1520_;
  wire _1521_;
  wire _1522_;
  wire _1523_;
  wire _1524_;
  wire _1525_;
  wire _1526_;
  wire _1527_;
  wire _1528_;
  wire _1529_;
  wire _1530_;
  wire _1531_;
  wire _1532_;
  wire _1533_;
  wire _1534_;
  wire _1535_;
  wire _1536_;
  wire _1537_;
  wire _1538_;
  wire _1539_;
  wire _1540_;
  wire _1541_;
  wire _1542_;
  wire _1543_;
  wire _1544_;
  wire _1545_;
  wire _1546_;
  wire _1547_;
  wire _1548_;
  wire _1549_;
  wire _1550_;
  wire _1551_;
  wire _1552_;
  wire _1553_;
  wire _1554_;
  wire _1555_;
  wire _1556_;
  wire _1557_;
  wire _1558_;
  wire _1559_;
  wire _1560_;
  wire _1561_;
  wire _1562_;
  wire _1563_;
  wire _1564_;
  wire _1565_;
  wire _1566_;
  wire _1567_;
  wire _1568_;
  wire _1569_;
  wire _1570_;
  wire _1571_;
  wire _1572_;
  wire _1573_;
  wire _1574_;
  wire _1575_;
  wire _1576_;
  wire _1577_;
  wire _1578_;
  wire _1579_;
  wire _1580_;
  wire _1581_;
  wire _1582_;
  wire _1583_;
  wire _1584_;
  wire _1585_;
  wire _1586_;
  wire _1587_;
  wire _1588_;
  wire _1589_;
  wire _1590_;
  wire _1591_;
  wire _1592_;
  wire _1593_;
  wire _1594_;
  wire _1595_;
  wire _1596_;
  wire _1597_;
  wire _1598_;
  wire _1599_;
  wire _1600_;
  wire _1601_;
  wire _1602_;
  wire _1603_;
  wire _1604_;
  wire _1605_;
  wire _1606_;
  wire _1607_;
  wire _1608_;
  wire _1609_;
  wire _1610_;
  wire _1611_;
  wire _1612_;
  wire _1613_;
  wire _1614_;
  wire _1615_;
  wire _1616_;
  wire _1617_;
  wire _1618_;
  wire _1619_;
  wire _1620_;
  wire _1621_;
  wire _1622_;
  wire _1623_;
  wire _1624_;
  wire _1625_;
  wire _1626_;
  wire _1627_;
  wire _1628_;
  wire _1629_;
  wire _1630_;
  wire _1631_;
  wire _1632_;
  wire _1633_;
  wire _1634_;
  wire _1635_;
  wire _1636_;
  wire _1637_;
  wire _1638_;
  wire _1639_;
  wire _1640_;
  wire _1641_;
  wire _1642_;
  wire _1643_;
  wire _1644_;
  wire _1645_;
  wire _1646_;
  wire _1647_;
  wire _1648_;
  wire _1649_;
  wire _1650_;
  wire _1651_;
  wire _1652_;
  wire _1653_;
  wire _1654_;
  wire _1655_;
  wire _1656_;
  wire _1657_;
  wire _1658_;
  wire _1659_;
  wire _1660_;
  wire _1661_;
  wire _1662_;
  wire _1663_;
  wire _1664_;
  wire _1665_;
  wire _1666_;
  wire _1667_;
  wire _1668_;
  wire _1669_;
  wire _1670_;
  wire _1671_;
  wire _1672_;
  wire _1673_;
  wire _1674_;
  wire _1675_;
  wire _1676_;
  wire _1677_;
  wire _1678_;
  wire _1679_;
  wire _1680_;
  wire _1681_;
  wire _1682_;
  wire _1683_;
  wire _1684_;
  wire _1685_;
  wire _1686_;
  wire _1687_;
  wire _1688_;
  wire _1689_;
  wire _1690_;
  wire _1691_;
  wire _1692_;
  wire _1693_;
  wire _1694_;
  wire _1695_;
  wire _1696_;
  wire _1697_;
  wire _1698_;
  wire _1699_;
  wire _1700_;
  wire _1701_;
  wire _1702_;
  wire _1703_;
  wire _1704_;
  wire _1705_;
  wire _1706_;
  wire _1707_;
  wire _1708_;
  wire _1709_;
  wire _1710_;
  wire _1711_;
  wire _1712_;
  wire _1713_;
  wire _1714_;
  wire _1715_;
  wire _1716_;
  wire _1717_;
  wire _1718_;
  wire _1719_;
  wire _1720_;
  wire _1721_;
  wire _1722_;
  wire _1723_;
  wire _1724_;
  wire _1725_;
  wire _1726_;
  wire _1727_;
  wire _1728_;
  wire _1729_;
  wire _1730_;
  wire _1731_;
  wire _1732_;
  wire _1733_;
  wire _1734_;
  wire _1735_;
  wire _1736_;
  wire _1737_;
  wire _1738_;
  wire _1739_;
  wire _1740_;
  wire _1741_;
  wire _1742_;
  wire _1743_;
  wire _1744_;
  wire _1745_;
  wire _1746_;
  wire _1747_;
  wire _1748_;
  wire _1749_;
  wire _1750_;
  wire _1751_;
  wire _1752_;
  wire _1753_;
  wire _1754_;
  wire _1755_;
  wire _1756_;
  wire _1757_;
  wire _1758_;
  wire _1759_;
  wire _1760_;
  wire _1761_;
  wire _1762_;
  wire _1763_;
  wire _1764_;
  wire _1765_;
  wire _1766_;
  wire _1767_;
  wire _1768_;
  wire _1769_;
  wire _1770_;
  wire _1771_;
  wire _1772_;
  wire _1773_;
  wire _1774_;
  wire _1775_;
  wire _1776_;
  wire _1777_;
  wire _1778_;
  wire _1779_;
  wire _1780_;
  wire _1781_;
  wire _1782_;
  wire _1783_;
  wire _1784_;
  wire _1785_;
  wire _1786_;
  wire _1787_;
  wire _1788_;
  wire _1789_;
  wire _1790_;
  wire _1791_;
  wire _1792_;
  wire _1793_;
  wire _1794_;
  wire _1795_;
  wire _1796_;
  wire _1797_;
  wire _1798_;
  wire _1799_;
  wire _1800_;
  wire _1801_;
  wire _1802_;
  wire _1803_;
  wire _1804_;
  wire _1805_;
  wire _1806_;
  wire _1807_;
  wire _1808_;
  wire _1809_;
  wire _1810_;
  wire _1811_;
  wire _1812_;
  wire _1813_;
  wire _1814_;
  wire _1815_;
  wire _1816_;
  wire _1817_;
  wire _1818_;
  wire _1819_;
  wire _1820_;
  wire _1821_;
  wire _1822_;
  wire _1823_;
  wire _1824_;
  wire _1825_;
  wire _1826_;
  wire _1827_;
  wire _1828_;
  wire _1829_;
  wire _1830_;
  wire _1831_;
  wire _1832_;
  wire _1833_;
  wire _1834_;
  wire _1835_;
  wire _1836_;
  wire _1837_;
  wire _1838_;
  wire _1839_;
  wire _1840_;
  wire _1841_;
  wire _1842_;
  wire _1843_;
  wire _1844_;
  wire _1845_;
  wire _1846_;
  wire _1847_;
  wire _1848_;
  wire _1849_;
  wire _1850_;
  wire _1851_;
  wire _1852_;
  wire _1853_;
  wire _1854_;
  wire _1855_;
  wire _1856_;
  wire _1857_;
  wire _1858_;
  wire _1859_;
  wire _1860_;
  wire _1861_;
  wire _1862_;
  wire _1863_;
  wire _1864_;
  wire _1865_;
  wire _1866_;
  wire _1867_;
  wire _1868_;
  wire _1869_;
  wire _1870_;
  wire _1871_;
  wire _1872_;
  wire _1873_;
  wire _1874_;
  wire _1875_;
  wire _1876_;
  wire _1877_;
  wire _1878_;
  wire _1879_;
  wire _1880_;
  wire _1881_;
  wire _1882_;
  wire _1883_;
  wire _1884_;
  wire _1885_;
  wire _1886_;
  wire _1887_;
  wire _1888_;
  wire _1889_;
  wire _1890_;
  wire _1891_;
  wire _1892_;
  wire _1893_;
  wire _1894_;
  wire _1895_;
  wire _1896_;
  wire _1897_;
  wire _1898_;
  wire _1899_;
  wire _1900_;
  wire _1901_;
  wire _1902_;
  wire _1903_;
  wire _1904_;
  wire _1905_;
  wire _1906_;
  wire _1907_;
  wire _1908_;
  wire _1909_;
  wire _1910_;
  wire _1911_;
  wire _1912_;
  wire _1913_;
  wire _1914_;
  wire _1915_;
  wire _1916_;
  wire _1917_;
  wire _1918_;
  wire _1919_;
  wire _1920_;
  wire _1921_;
  wire _1922_;
  wire _1923_;
  wire _1924_;
  wire _1925_;
  wire _1926_;
  wire _1927_;
  wire _1928_;
  wire _1929_;
  wire _1930_;
  wire _1931_;
  wire _1932_;
  wire _1933_;
  wire _1934_;
  wire _1935_;
  wire _1936_;
  wire _1937_;
  wire _1938_;
  wire _1939_;
  wire _1940_;
  wire _1941_;
  wire _1942_;
  wire _1943_;
  wire _1944_;
  wire _1945_;
  wire _1946_;
  wire _1947_;
  wire _1948_;
  wire _1949_;
  wire _1950_;
  wire _1951_;
  wire _1952_;
  wire _1953_;
  wire _1954_;
  wire _1955_;
  wire _1956_;
  wire _1957_;
  wire _1958_;
  wire _1959_;
  wire _1960_;
  wire _1961_;
  wire _1962_;
  wire _1963_;
  wire _1964_;
  wire _1965_;
  wire _1966_;
  wire _1967_;
  wire _1968_;
  wire _1969_;
  wire _1970_;
  wire _1971_;
  wire _1972_;
  wire _1973_;
  wire _1974_;
  wire _1975_;
  wire _1976_;
  wire _1977_;
  wire _1978_;
  wire _1979_;
  wire _1980_;
  wire _1981_;
  wire _1982_;
  wire _1983_;
  wire _1984_;
  wire _1985_;
  wire _1986_;
  wire _1987_;
  wire _1988_;
  wire _1989_;
  wire _1990_;
  wire _1991_;
  wire _1992_;
  wire _1993_;
  wire _1994_;
  wire _1995_;
  wire _1996_;
  wire _1997_;
  wire _1998_;
  wire _1999_;
  wire _2000_;
  wire _2001_;
  wire _2002_;
  wire _2003_;
  wire _2004_;
  wire _2005_;
  wire _2006_;
  wire _2007_;
  wire _2008_;
  wire _2009_;
  wire _2010_;
  wire _2011_;
  wire _2012_;
  wire _2013_;
  wire _2014_;
  wire _2015_;
  wire _2016_;
  wire _2017_;
  wire _2018_;
  wire _2019_;
  wire _2020_;
  wire _2021_;
  wire _2022_;
  wire _2023_;
  wire _2024_;
  wire _2025_;
  wire _2026_;
  wire _2027_;
  wire _2028_;
  wire _2029_;
  wire _2030_;
  wire _2031_;
  wire _2032_;
  wire _2033_;
  wire _2034_;
  wire _2035_;
  wire _2036_;
  wire _2037_;
  wire _2038_;
  wire _2039_;
  wire _2040_;
  wire _2041_;
  wire _2042_;
  wire _2043_;
  wire _2044_;
  wire _2045_;
  wire _2046_;
  wire _2047_;
  wire _2048_;
  wire _2049_;
  wire _2050_;
  wire _2051_;
  wire _2052_;
  wire _2053_;
  wire _2054_;
  wire _2055_;
  wire _2056_;
  wire _2057_;
  wire _2058_;
  wire _2059_;
  wire _2060_;
  wire _2061_;
  wire _2062_;
  wire _2063_;
  wire _2064_;
  wire _2065_;
  wire _2066_;
  wire _2067_;
  wire _2068_;
  wire _2069_;
  wire _2070_;
  wire _2071_;
  wire _2072_;
  wire _2073_;
  wire _2074_;
  wire _2075_;
  wire _2076_;
  wire _2077_;
  wire _2078_;
  wire _2079_;
  wire _2080_;
  wire _2081_;
  wire _2082_;
  wire _2083_;
  wire _2084_;
  wire _2085_;
  wire _2086_;
  wire _2087_;
  wire _2088_;
  wire _2089_;
  wire _2090_;
  wire _2091_;
  wire _2092_;
  wire _2093_;
  wire _2094_;
  wire _2095_;
  wire _2096_;
  wire _2097_;
  wire _2098_;
  wire _2099_;
  wire _2100_;
  wire _2101_;
  wire _2102_;
  wire _2103_;
  wire _2104_;
  wire _2105_;
  wire _2106_;
  wire _2107_;
  wire _2108_;
  wire _2109_;
  wire _2110_;
  wire _2111_;
  wire _2112_;
  wire _2113_;
  wire _2114_;
  wire _2115_;
  wire _2116_;
  wire _2117_;
  wire _2118_;
  wire _2119_;
  wire _2120_;
  wire _2121_;
  wire _2122_;
  wire _2123_;
  wire _2124_;
  wire _2125_;
  wire _2126_;
  wire _2127_;
  wire _2128_;
  wire _2129_;
  wire _2130_;
  wire _2131_;
  wire _2132_;
  wire _2133_;
  wire _2134_;
  wire _2135_;
  wire _2136_;
  wire _2137_;
  wire _2138_;
  wire _2139_;
  wire _2140_;
  wire _2141_;
  wire _2142_;
  wire _2143_;
  wire _2144_;
  wire _2145_;
  wire _2146_;
  wire _2147_;
  wire _2148_;
  wire _2149_;
  wire _2150_;
  wire _2151_;
  wire _2152_;
  wire _2153_;
  wire _2154_;
  wire _2155_;
  wire _2156_;
  wire _2157_;
  wire _2158_;
  wire _2159_;
  wire _2160_;
  wire _2161_;
  wire _2162_;
  wire _2163_;
  wire _2164_;
  wire _2165_;
  wire _2166_;
  wire _2167_;
  wire _2168_;
  wire _2169_;
  wire _2170_;
  wire _2171_;
  wire _2172_;
  wire _2173_;
  wire _2174_;
  wire _2175_;
  wire _2176_;
  wire _2177_;
  wire _2178_;
  wire _2179_;
  wire _2180_;
  wire _2181_;
  wire _2182_;
  wire _2183_;
  wire _2184_;
  wire _2185_;
  wire _2186_;
  wire _2187_;
  wire _2188_;
  wire _2189_;
  wire _2190_;
  wire _2191_;
  wire _2192_;
  wire _2193_;
  wire _2194_;
  wire _2195_;
  wire _2196_;
  wire _2197_;
  wire _2198_;
  wire _2199_;
  wire _2200_;
  wire _2201_;
  wire _2202_;
  wire _2203_;
  wire _2204_;
  wire _2205_;
  wire _2206_;
  wire _2207_;
  wire _2208_;
  wire _2209_;
  wire _2210_;
  wire _2211_;
  wire _2212_;
  wire _2213_;
  wire _2214_;
  wire _2215_;
  wire _2216_;
  wire _2217_;
  wire _2218_;
  wire _2219_;
  wire _2220_;
  wire _2221_;
  wire _2222_;
  wire _2223_;
  wire _2224_;
  wire _2225_;
  wire _2226_;
  wire _2227_;
  wire _2228_;
  wire _2229_;
  wire _2230_;
  wire _2231_;
  wire _2232_;
  wire _2233_;
  wire _2234_;
  wire _2235_;
  wire _2236_;
  wire _2237_;
  wire _2238_;
  wire _2239_;
  wire _2240_;
  wire _2241_;
  wire _2242_;
  wire _2243_;
  wire _2244_;
  wire _2245_;
  wire _2246_;
  wire _2247_;
  wire _2248_;
  wire _2249_;
  wire _2250_;
  wire _2251_;
  wire _2252_;
  wire _2253_;
  wire _2254_;
  wire _2255_;
  wire _2256_;
  wire _2257_;
  wire _2258_;
  wire _2259_;
  wire _2260_;
  wire _2261_;
  wire _2262_;
  wire _2263_;
  wire _2264_;
  wire _2265_;
  wire _2266_;
  wire _2267_;
  wire _2268_;
  wire _2269_;
  wire _2270_;
  wire _2271_;
  wire _2272_;
  wire _2273_;
  wire _2274_;
  wire _2275_;
  wire _2276_;
  wire _2277_;
  wire _2278_;
  wire _2279_;
  wire _2280_;
  wire _2281_;
  wire _2282_;
  wire _2283_;
  wire _2284_;
  wire _2285_;
  wire _2286_;
  wire _2287_;
  wire _2288_;
  wire _2289_;
  wire _2290_;
  wire _2291_;
  wire _2292_;
  wire _2293_;
  wire _2294_;
  wire _2295_;
  wire _2296_;
  wire _2297_;
  wire _2298_;
  wire _2299_;
  wire _2300_;
  wire _2301_;
  wire _2302_;
  wire _2303_;
  wire _2304_;
  wire _2305_;
  wire _2306_;
  wire _2307_;
  wire _2308_;
  wire _2309_;
  wire _2310_;
  wire _2311_;
  wire _2312_;
  wire _2313_;
  wire _2314_;
  wire _2315_;
  wire _2316_;
  wire _2317_;
  wire _2318_;
  wire _2319_;
  wire _2320_;
  wire _2321_;
  wire _2322_;
  wire _2323_;
  wire _2324_;
  wire _2325_;
  wire _2326_;
  wire _2327_;
  wire _2328_;
  wire _2329_;
  wire _2330_;
  wire _2331_;
  wire _2332_;
  wire _2333_;
  wire _2334_;
  wire _2335_;
  wire _2336_;
  wire _2337_;
  wire _2338_;
  wire _2339_;
  wire _2340_;
  wire _2341_;
  wire _2342_;
  wire _2343_;
  wire _2344_;
  wire _2345_;
  wire _2346_;
  wire _2347_;
  wire _2348_;
  wire _2349_;
  wire _2350_;
  wire _2351_;
  wire _2352_;
  wire _2353_;
  wire _2354_;
  wire _2355_;
  wire _2356_;
  wire _2357_;
  wire _2358_;
  wire _2359_;
  wire _2360_;
  wire _2361_;
  wire _2362_;
  wire _2363_;
  wire _2364_;
  wire _2365_;
  wire _2366_;
  wire _2367_;
  wire _2368_;
  wire _2369_;
  wire _2370_;
  wire _2371_;
  wire _2372_;
  wire _2373_;
  wire _2374_;
  wire _2375_;
  wire _2376_;
  wire _2377_;
  wire _2378_;
  wire _2379_;
  wire _2380_;
  wire _2381_;
  wire _2382_;
  wire _2383_;
  wire _2384_;
  wire _2385_;
  wire _2386_;
  wire _2387_;
  wire _2388_;
  wire _2389_;
  wire _2390_;
  wire _2391_;
  wire _2392_;
  wire _2393_;
  wire _2394_;
  wire _2395_;
  wire _2396_;
  wire _2397_;
  wire _2398_;
  wire _2399_;
  wire _2400_;
  wire _2401_;
  wire _2402_;
  wire _2403_;
  wire _2404_;
  wire _2405_;
  wire _2406_;
  wire _2407_;
  wire _2408_;
  wire _2409_;
  wire _2410_;
  wire _2411_;
  wire _2412_;
  wire _2413_;
  wire _2414_;
  wire _2415_;
  wire _2416_;
  wire _2417_;
  wire _2418_;
  wire _2419_;
  wire _2420_;
  wire _2421_;
  wire _2422_;
  wire _2423_;
  wire _2424_;
  wire _2425_;
  wire _2426_;
  wire _2427_;
  wire _2428_;
  wire _2429_;
  wire _2430_;
  wire _2431_;
  wire _2432_;
  wire _2433_;
  wire _2434_;
  wire _2435_;
  wire _2436_;
  wire _2437_;
  wire _2438_;
  wire _2439_;
  wire _2440_;
  wire _2441_;
  wire _2442_;
  wire _2443_;
  wire _2444_;
  wire _2445_;
  wire _2446_;
  wire _2447_;
  wire _2448_;
  wire _2449_;
  wire _2450_;
  wire _2451_;
  wire _2452_;
  wire _2453_;
  wire _2454_;
  wire _2455_;
  wire _2456_;
  wire _2457_;
  wire _2458_;
  wire _2459_;
  wire _2460_;
  wire _2461_;
  wire _2462_;
  wire _2463_;
  wire _2464_;
  wire _2465_;
  wire _2466_;
  wire _2467_;
  wire _2468_;
  wire _2469_;
  wire _2470_;
  wire _2471_;
  wire _2472_;
  wire _2473_;
  wire _2474_;
  wire _2475_;
  wire _2476_;
  wire _2477_;
  wire _2478_;
  wire _2479_;
  wire _2480_;
  wire _2481_;
  wire _2482_;
  wire _2483_;
  wire _2484_;
  wire _2485_;
  wire _2486_;
  wire _2487_;
  wire _2488_;
  wire _2489_;
  wire _2490_;
  wire _2491_;
  wire _2492_;
  wire _2493_;
  wire _2494_;
  wire _2495_;
  wire _2496_;
  wire _2497_;
  wire _2498_;
  wire _2499_;
  wire _2500_;
  wire _2501_;
  wire _2502_;
  wire _2503_;
  wire _2504_;
  wire _2505_;
  wire _2506_;
  wire _2507_;
  wire _2508_;
  wire _2509_;
  wire _2510_;
  wire _2511_;
  wire _2512_;
  wire _2513_;
  wire _2514_;
  wire _2515_;
  wire _2516_;
  wire _2517_;
  wire _2518_;
  wire _2519_;
  wire _2520_;
  wire _2521_;
  wire _2522_;
  wire _2523_;
  wire _2524_;
  wire _2525_;
  wire _2526_;
  wire _2527_;
  wire _2528_;
  wire _2529_;
  wire _2530_;
  wire _2531_;
  wire _2532_;
  wire _2533_;
  wire _2534_;
  wire _2535_;
  wire _2536_;
  wire _2537_;
  wire _2538_;
  wire _2539_;
  wire _2540_;
  wire _2541_;
  wire _2542_;
  wire _2543_;
  wire _2544_;
  wire _2545_;
  wire _2546_;
  wire _2547_;
  wire _2548_;
  wire _2549_;
  wire _2550_;
  wire _2551_;
  wire _2552_;
  wire _2553_;
  wire _2554_;
  wire _2555_;
  wire _2556_;
  wire _2557_;
  wire _2558_;
  wire _2559_;
  wire _2560_;
  wire _2561_;
  wire _2562_;
  wire _2563_;
  wire _2564_;
  wire _2565_;
  wire _2566_;
  wire _2567_;
  wire _2568_;
  wire _2569_;
  wire _2570_;
  wire _2571_;
  wire _2572_;
  wire _2573_;
  wire _2574_;
  wire _2575_;
  wire _2576_;
  wire _2577_;
  wire _2578_;
  wire _2579_;
  wire _2580_;
  wire _2581_;
  wire _2582_;
  wire _2583_;
  wire _2584_;
  wire _2585_;
  wire _2586_;
  wire _2587_;
  wire _2588_;
  wire _2589_;
  wire _2590_;
  wire _2591_;
  wire _2592_;
  wire _2593_;
  wire _2594_;
  wire _2595_;
  wire _2596_;
  wire _2597_;
  wire _2598_;
  wire _2599_;
  wire _2600_;
  wire _2601_;
  wire _2602_;
  wire _2603_;
  wire _2604_;
  wire _2605_;
  wire _2606_;
  wire _2607_;
  wire _2608_;
  wire _2609_;
  wire _2610_;
  wire _2611_;
  wire _2612_;
  wire _2613_;
  wire _2614_;
  wire _2615_;
  wire _2616_;
  wire _2617_;
  wire _2618_;
  wire _2619_;
  wire _2620_;
  wire _2621_;
  wire _2622_;
  wire _2623_;
  wire _2624_;
  wire _2625_;
  wire _2626_;
  wire _2627_;
  wire _2628_;
  wire _2629_;
  wire _2630_;
  wire _2631_;
  wire _2632_;
  wire _2633_;
  wire _2634_;
  wire _2635_;
  wire _2636_;
  wire _2637_;
  wire _2638_;
  wire _2639_;
  wire _2640_;
  wire _2641_;
  wire _2642_;
  wire _2643_;
  wire _2644_;
  wire _2645_;
  wire _2646_;
  wire _2647_;
  wire _2648_;
  wire _2649_;
  wire _2650_;
  wire _2651_;
  wire _2652_;
  wire _2653_;
  wire _2654_;
  wire _2655_;
  wire _2656_;
  wire _2657_;
  wire _2658_;
  wire _2659_;
  wire _2660_;
  wire _2661_;
  wire _2662_;
  wire _2663_;
  wire _2664_;
  wire _2665_;
  wire _2666_;
  wire _2667_;
  wire _2668_;
  wire _2669_;
  wire _2670_;
  wire _2671_;
  wire _2672_;
  wire _2673_;
  wire _2674_;
  wire _2675_;
  wire _2676_;
  wire _2677_;
  wire _2678_;
  wire _2679_;
  wire _2680_;
  wire _2681_;
  wire _2682_;
  wire _2683_;
  wire _2684_;
  wire _2685_;
  wire _2686_;
  wire _2687_;
  wire _2688_;
  wire _2689_;
  wire _2690_;
  wire _2691_;
  wire _2692_;
  wire _2693_;
  wire _2694_;
  wire _2695_;
  wire _2696_;
  wire _2697_;
  wire _2698_;
  wire _2699_;
  wire _2700_;
  wire _2701_;
  wire _2702_;
  wire _2703_;
  wire _2704_;
  wire _2705_;
  wire _2706_;
  wire _2707_;
  wire _2708_;
  wire _2709_;
  wire _2710_;
  wire _2711_;
  wire _2712_;
  wire _2713_;
  wire _2714_;
  wire _2715_;
  wire _2716_;
  wire _2717_;
  wire _2718_;
  wire _2719_;
  wire _2720_;
  wire _2721_;
  wire _2722_;
  wire _2723_;
  wire _2724_;
  wire _2725_;
  wire _2726_;
  wire _2727_;
  wire _2728_;
  wire _2729_;
  wire _2730_;
  wire _2731_;
  wire _2732_;
  wire _2733_;
  wire _2734_;
  wire _2735_;
  wire _2736_;
  wire _2737_;
  wire _2738_;
  wire _2739_;
  wire _2740_;
  wire _2741_;
  wire _2742_;
  wire _2743_;
  wire _2744_;
  wire _2745_;
  wire _2746_;
  wire _2747_;
  wire _2748_;
  wire _2749_;
  wire _2750_;
  wire _2751_;
  wire _2752_;
  wire _2753_;
  wire _2754_;
  wire _2755_;
  wire _2756_;
  wire _2757_;
  wire _2758_;
  wire _2759_;
  wire _2760_;
  wire _2761_;
  wire _2762_;
  wire _2763_;
  wire _2764_;
  wire _2765_;
  wire _2766_;
  wire _2767_;
  wire _2768_;
  wire _2769_;
  wire _2770_;
  wire _2771_;
  wire _2772_;
  wire _2773_;
  wire _2774_;
  wire _2775_;
  wire _2776_;
  wire _2777_;
  wire _2778_;
  wire _2779_;
  wire _2780_;
  wire _2781_;
  wire _2782_;
  wire _2783_;
  wire _2784_;
  wire _2785_;
  wire _2786_;
  wire _2787_;
  wire _2788_;
  wire _2789_;
  wire _2790_;
  wire _2791_;
  wire _2792_;
  wire _2793_;
  wire _2794_;
  wire _2795_;
  wire _2796_;
  wire _2797_;
  wire _2798_;
  wire _2799_;
  wire _2800_;
  wire _2801_;
  wire _2802_;
  wire _2803_;
  wire _2804_;
  wire _2805_;
  wire _2806_;
  wire _2807_;
  wire _2808_;
  wire _2809_;
  wire _2810_;
  wire _2811_;
  wire _2812_;
  wire _2813_;
  wire _2814_;
  wire _2815_;
  wire _2816_;
  wire _2817_;
  wire _2818_;
  wire _2819_;
  wire _2820_;
  wire _2821_;
  wire _2822_;
  wire _2823_;
  wire _2824_;
  wire _2825_;
  wire _2826_;
  wire _2827_;
  wire _2828_;
  wire _2829_;
  wire _2830_;
  wire _2831_;
  wire _2832_;
  wire _2833_;
  wire _2834_;
  wire _2835_;
  wire _2836_;
  wire _2837_;
  wire _2838_;
  wire _2839_;
  wire _2840_;
  wire _2841_;
  wire _2842_;
  wire _2843_;
  wire _2844_;
  wire _2845_;
  wire _2846_;
  wire _2847_;
  wire _2848_;
  wire _2849_;
  wire _2850_;
  wire _2851_;
  wire _2852_;
  wire _2853_;
  wire _2854_;
  wire _2855_;
  wire _2856_;
  wire _2857_;
  wire _2858_;
  wire _2859_;
  wire _2860_;
  wire _2861_;
  wire _2862_;
  wire _2863_;
  wire _2864_;
  wire _2865_;
  wire _2866_;
  wire _2867_;
  wire _2868_;
  wire _2869_;
  wire _2870_;
  wire _2871_;
  wire _2872_;
  wire _2873_;
  wire _2874_;
  wire _2875_;
  wire _2876_;
  wire _2877_;
  wire _2878_;
  wire _2879_;
  wire _2880_;
  wire _2881_;
  wire _2882_;
  wire _2883_;
  wire _2884_;
  wire _2885_;
  wire _2886_;
  wire _2887_;
  wire _2888_;
  wire _2889_;
  wire _2890_;
  wire _2891_;
  wire _2892_;
  wire _2893_;
  wire _2894_;
  wire _2895_;
  wire _2896_;
  wire _2897_;
  wire _2898_;
  wire _2899_;
  wire _2900_;
  wire _2901_;
  wire _2902_;
  wire _2903_;
  wire _2904_;
  wire _2905_;
  wire _2906_;
  wire _2907_;
  wire _2908_;
  wire _2909_;
  wire _2910_;
  wire _2911_;
  wire _2912_;
  wire _2913_;
  wire _2914_;
  wire _2915_;
  wire _2916_;
  wire _2917_;
  wire _2918_;
  wire _2919_;
  wire _2920_;
  wire _2921_;
  wire _2922_;
  wire _2923_;
  wire _2924_;
  wire _2925_;
  wire _2926_;
  wire _2927_;
  wire _2928_;
  wire _2929_;
  wire _2930_;
  wire _2931_;
  wire _2932_;
  wire _2933_;
  wire _2934_;
  wire _2935_;
  wire _2936_;
  wire _2937_;
  wire _2938_;
  wire _2939_;
  wire _2940_;
  wire _2941_;
  wire _2942_;
  wire _2943_;
  wire _2944_;
  wire _2945_;
  wire _2946_;
  wire _2947_;
  wire _2948_;
  wire _2949_;
  wire _2950_;
  wire _2951_;
  wire _2952_;
  wire _2953_;
  wire _2954_;
  wire _2955_;
  wire _2956_;
  wire _2957_;
  wire _2958_;
  wire _2959_;
  wire _2960_;
  wire _2961_;
  wire _2962_;
  wire _2963_;
  wire _2964_;
  wire _2965_;
  wire _2966_;
  wire _2967_;
  wire _2968_;
  wire _2969_;
  wire _2970_;
  wire _2971_;
  wire _2972_;
  wire _2973_;
  wire _2974_;
  wire _2975_;
  wire _2976_;
  wire _2977_;
  wire _2978_;
  wire _2979_;
  wire _2980_;
  wire _2981_;
  wire _2982_;
  wire _2983_;
  wire _2984_;
  wire _2985_;
  wire _2986_;
  input [127:0] cipher_key;
  wire [127:0] cipher_key;
  output [127:0] ciphertext;
  wire [127:0] ciphertext;
  input clk;
  wire clk;
  output encrypt_done;
  wire encrypt_done;
  input encrypt_start;
  wire encrypt_start;
  wire encrypting;
  input [127:0] plaintext;
  wire [127:0] plaintext;
  wire [2:0] round_counter;
  wire [127:0] round_key;
  input rst;
  wire rst;
  wire [127:0] state;
    not _2987_(_0001_, rst);
    and _2988_(_0778_, round_counter[1], round_counter[0]);
    nand _2989_(_0779_, _0778_, round_counter[2]);
    not _2990_(_0780_, encrypting);
    nand _2991_(_0781_, encrypt_start, _0780_);
    and _2992_(_0782_, _0781_, encrypting);
    and _2993_(_0783_, _0782_, _0779_);
    and _2994_(_0784_, _0783_, encrypt_done);
    and _2995_(_0785_, _0778_, round_counter[2]);
    and _2996_(_0786_, _0785_, encrypting);
    and _2997_(_0787_, _0786_, _0781_);
    not _2998_(_0788_, _0787_);
    nor _2999_(_0789_, _0788_, _0783_);
    or _3000_(_0390_, _0789_, _0784_);
    or _3001_(_0790_, encrypt_start, encrypting);
    nand _3002_(_0791_, _0782_, _0785_);
    nand _3003_(_0792_, _0791_, _0790_);
    and _3004_(_0793_, _0792_, state[0]);
    and _3005_(_0794_, _0791_, _0790_);
    xor _3006_(_0795_, round_key[0], state[0]);
    and _3007_(_0796_, _0795_, _0779_);
    and _3008_(_0797_, _0796_, encrypting);
    and _3009_(_0798_, _0797_, _0781_);
    not _3010_(_0799_, _0781_);
    and _3011_(_0800_, _0799_, plaintext[0]);
    or _3012_(_0801_, _0800_, _0798_);
    and _3013_(_0802_, _0801_, _0794_);
    or _3014_(_0391_, _0802_, _0793_);
    and _3015_(_0803_, _0792_, state[1]);
    xor _3016_(_0804_, round_key[1], state[1]);
    and _3017_(_0805_, _0804_, _0779_);
    and _3018_(_0806_, _0805_, encrypting);
    and _3019_(_0807_, _0806_, _0781_);
    and _3020_(_0808_, _0799_, plaintext[1]);
    or _3021_(_0809_, _0808_, _0807_);
    and _3022_(_0810_, _0809_, _0794_);
    or _3023_(_0392_, _0810_, _0803_);
    and _3024_(_0811_, _0792_, state[2]);
    xor _3025_(_0812_, round_key[2], state[2]);
    and _3026_(_0813_, _0812_, _0779_);
    and _3027_(_0814_, _0813_, encrypting);
    and _3028_(_0815_, _0814_, _0781_);
    and _3029_(_0816_, _0799_, plaintext[2]);
    or _3030_(_0817_, _0816_, _0815_);
    and _3031_(_0818_, _0817_, _0794_);
    or _3032_(_0393_, _0818_, _0811_);
    and _3033_(_0819_, _0792_, state[3]);
    xor _3034_(_0820_, round_key[3], state[3]);
    and _3035_(_0821_, _0820_, _0779_);
    and _3036_(_0822_, _0821_, encrypting);
    and _3037_(_0823_, _0822_, _0781_);
    and _3038_(_0824_, _0799_, plaintext[3]);
    or _3039_(_0825_, _0824_, _0823_);
    and _3040_(_0826_, _0825_, _0794_);
    or _3041_(_0394_, _0826_, _0819_);
    and _3042_(_0827_, _0792_, state[4]);
    xor _3043_(_0828_, round_key[4], state[4]);
    and _3044_(_0829_, _0828_, _0779_);
    and _3045_(_0830_, _0829_, encrypting);
    and _3046_(_0831_, _0830_, _0781_);
    and _3047_(_0832_, _0799_, plaintext[4]);
    or _3048_(_0833_, _0832_, _0831_);
    and _3049_(_0834_, _0833_, _0794_);
    or _3050_(_0395_, _0834_, _0827_);
    and _3051_(_0835_, _0792_, state[5]);
    xor _3052_(_0836_, round_key[5], state[5]);
    and _3053_(_0837_, _0836_, _0779_);
    and _3054_(_0838_, _0837_, encrypting);
    and _3055_(_0839_, _0838_, _0781_);
    and _3056_(_0840_, _0799_, plaintext[5]);
    or _3057_(_0841_, _0840_, _0839_);
    and _3058_(_0842_, _0841_, _0794_);
    or _3059_(_0396_, _0842_, _0835_);
    and _3060_(_0843_, _0792_, state[6]);
    xor _3061_(_0844_, round_key[6], state[6]);
    and _3062_(_0845_, _0844_, _0779_);
    and _3063_(_0846_, _0845_, encrypting);
    and _3064_(_0847_, _0846_, _0781_);
    and _3065_(_0848_, _0799_, plaintext[6]);
    or _3066_(_0849_, _0848_, _0847_);
    and _3067_(_0850_, _0849_, _0794_);
    or _3068_(_0397_, _0850_, _0843_);
    and _3069_(_0851_, _0792_, state[7]);
    xor _3070_(_0852_, round_key[7], state[7]);
    and _3071_(_0853_, _0852_, _0779_);
    and _3072_(_0854_, _0853_, encrypting);
    and _3073_(_0855_, _0854_, _0781_);
    and _3074_(_0856_, _0799_, plaintext[7]);
    or _3075_(_0857_, _0856_, _0855_);
    and _3076_(_0858_, _0857_, _0794_);
    or _3077_(_0398_, _0858_, _0851_);
    and _3078_(_0859_, _0792_, state[8]);
    xor _3079_(_0860_, round_key[8], state[8]);
    and _3080_(_0861_, _0860_, _0779_);
    and _3081_(_0862_, _0861_, encrypting);
    and _3082_(_0863_, _0862_, _0781_);
    and _3083_(_0864_, _0799_, plaintext[8]);
    or _3084_(_0865_, _0864_, _0863_);
    and _3085_(_0866_, _0865_, _0794_);
    or _3086_(_0399_, _0866_, _0859_);
    and _3087_(_0867_, _0792_, state[9]);
    xor _3088_(_0868_, round_key[9], state[9]);
    and _3089_(_0869_, _0868_, _0779_);
    and _3090_(_0870_, _0869_, encrypting);
    and _3091_(_0871_, _0870_, _0781_);
    and _3092_(_0872_, _0799_, plaintext[9]);
    or _3093_(_0873_, _0872_, _0871_);
    and _3094_(_0874_, _0873_, _0794_);
    or _3095_(_0400_, _0874_, _0867_);
    and _3096_(_0875_, _0792_, state[10]);
    xor _3097_(_0876_, round_key[10], state[10]);
    and _3098_(_0877_, _0876_, _0779_);
    and _3099_(_0878_, _0877_, encrypting);
    and _3100_(_0879_, _0878_, _0781_);
    and _3101_(_0880_, _0799_, plaintext[10]);
    or _3102_(_0881_, _0880_, _0879_);
    and _3103_(_0882_, _0881_, _0794_);
    or _3104_(_0401_, _0882_, _0875_);
    and _3105_(_0883_, _0792_, state[11]);
    xor _3106_(_0884_, round_key[11], state[11]);
    and _3107_(_0885_, _0884_, _0779_);
    and _3108_(_0886_, _0885_, encrypting);
    and _3109_(_0887_, _0886_, _0781_);
    and _3110_(_0888_, _0799_, plaintext[11]);
    or _3111_(_0889_, _0888_, _0887_);
    and _3112_(_0890_, _0889_, _0794_);
    or _3113_(_0402_, _0890_, _0883_);
    and _3114_(_0891_, _0792_, state[12]);
    xor _3115_(_0892_, round_key[12], state[12]);
    and _3116_(_0893_, _0892_, _0779_);
    and _3117_(_0894_, _0893_, encrypting);
    and _3118_(_0895_, _0894_, _0781_);
    and _3119_(_0896_, _0799_, plaintext[12]);
    or _3120_(_0897_, _0896_, _0895_);
    and _3121_(_0898_, _0897_, _0794_);
    or _3122_(_0403_, _0898_, _0891_);
    and _3123_(_0899_, _0792_, state[13]);
    xor _3124_(_0900_, round_key[13], state[13]);
    and _3125_(_0901_, _0900_, _0779_);
    and _3126_(_0902_, _0901_, encrypting);
    and _3127_(_0903_, _0902_, _0781_);
    and _3128_(_0904_, _0799_, plaintext[13]);
    or _3129_(_0905_, _0904_, _0903_);
    and _3130_(_0906_, _0905_, _0794_);
    or _3131_(_0404_, _0906_, _0899_);
    and _3132_(_0907_, _0792_, state[14]);
    xor _3133_(_0908_, round_key[14], state[14]);
    and _3134_(_0909_, _0908_, _0779_);
    and _3135_(_0910_, _0909_, encrypting);
    and _3136_(_0911_, _0910_, _0781_);
    and _3137_(_0912_, _0799_, plaintext[14]);
    or _3138_(_0913_, _0912_, _0911_);
    and _3139_(_0914_, _0913_, _0794_);
    or _3140_(_0405_, _0914_, _0907_);
    and _3141_(_0915_, _0792_, state[15]);
    xor _3142_(_0916_, round_key[15], state[15]);
    and _3143_(_0917_, _0916_, _0779_);
    and _3144_(_0918_, _0917_, encrypting);
    and _3145_(_0919_, _0918_, _0781_);
    and _3146_(_0920_, _0799_, plaintext[15]);
    or _3147_(_0921_, _0920_, _0919_);
    and _3148_(_0922_, _0921_, _0794_);
    or _3149_(_0406_, _0922_, _0915_);
    and _3150_(_0923_, _0792_, state[16]);
    xor _3151_(_0924_, round_key[16], state[16]);
    and _3152_(_0925_, _0924_, _0779_);
    and _3153_(_0926_, _0925_, encrypting);
    and _3154_(_0927_, _0926_, _0781_);
    and _3155_(_0928_, _0799_, plaintext[16]);
    or _3156_(_0929_, _0928_, _0927_);
    and _3157_(_0930_, _0929_, _0794_);
    or _3158_(_0407_, _0930_, _0923_);
    and _3159_(_0931_, _0792_, state[17]);
    xor _3160_(_0932_, round_key[17], state[17]);
    and _3161_(_0933_, _0932_, _0779_);
    and _3162_(_0934_, _0933_, encrypting);
    and _3163_(_0935_, _0934_, _0781_);
    and _3164_(_0936_, _0799_, plaintext[17]);
    or _3165_(_0937_, _0936_, _0935_);
    and _3166_(_0938_, _0937_, _0794_);
    or _3167_(_0408_, _0938_, _0931_);
    and _3168_(_0939_, _0792_, state[18]);
    xor _3169_(_0940_, round_key[18], state[18]);
    and _3170_(_0941_, _0940_, _0779_);
    and _3171_(_0942_, _0941_, encrypting);
    and _3172_(_0943_, _0942_, _0781_);
    and _3173_(_0944_, _0799_, plaintext[18]);
    or _3174_(_0945_, _0944_, _0943_);
    and _3175_(_0946_, _0945_, _0794_);
    or _3176_(_0409_, _0946_, _0939_);
    and _3177_(_0947_, _0792_, state[19]);
    xor _3178_(_0948_, round_key[19], state[19]);
    and _3179_(_0949_, _0948_, _0779_);
    and _3180_(_0950_, _0949_, encrypting);
    and _3181_(_0951_, _0950_, _0781_);
    and _3182_(_0952_, _0799_, plaintext[19]);
    or _3183_(_0953_, _0952_, _0951_);
    and _3184_(_0954_, _0953_, _0794_);
    or _3185_(_0410_, _0954_, _0947_);
    and _3186_(_0955_, _0792_, state[20]);
    xor _3187_(_0956_, round_key[20], state[20]);
    and _3188_(_0957_, _0956_, _0779_);
    and _3189_(_0958_, _0957_, encrypting);
    and _3190_(_0959_, _0958_, _0781_);
    and _3191_(_0960_, _0799_, plaintext[20]);
    or _3192_(_0961_, _0960_, _0959_);
    and _3193_(_0962_, _0961_, _0794_);
    or _3194_(_0411_, _0962_, _0955_);
    and _3195_(_0963_, _0792_, state[21]);
    xor _3196_(_0964_, round_key[21], state[21]);
    and _3197_(_0965_, _0964_, _0779_);
    and _3198_(_0966_, _0965_, encrypting);
    and _3199_(_0967_, _0966_, _0781_);
    and _3200_(_0968_, _0799_, plaintext[21]);
    or _3201_(_0969_, _0968_, _0967_);
    and _3202_(_0970_, _0969_, _0794_);
    or _3203_(_0412_, _0970_, _0963_);
    and _3204_(_0971_, _0792_, state[22]);
    xor _3205_(_0972_, round_key[22], state[22]);
    and _3206_(_0973_, _0972_, _0779_);
    and _3207_(_0974_, _0973_, encrypting);
    and _3208_(_0975_, _0974_, _0781_);
    and _3209_(_0976_, _0799_, plaintext[22]);
    or _3210_(_0977_, _0976_, _0975_);
    and _3211_(_0978_, _0977_, _0794_);
    or _3212_(_0413_, _0978_, _0971_);
    and _3213_(_0979_, _0792_, state[23]);
    xor _3214_(_0980_, round_key[23], state[23]);
    and _3215_(_0981_, _0980_, _0779_);
    and _3216_(_0982_, _0981_, encrypting);
    and _3217_(_0983_, _0982_, _0781_);
    and _3218_(_0984_, _0799_, plaintext[23]);
    or _3219_(_0985_, _0984_, _0983_);
    and _3220_(_0986_, _0985_, _0794_);
    or _3221_(_0414_, _0986_, _0979_);
    and _3222_(_0987_, _0792_, state[24]);
    xor _3223_(_0988_, round_key[24], state[24]);
    and _3224_(_0989_, _0988_, _0779_);
    and _3225_(_0990_, _0989_, encrypting);
    and _3226_(_0991_, _0990_, _0781_);
    and _3227_(_0992_, _0799_, plaintext[24]);
    or _3228_(_0993_, _0992_, _0991_);
    and _3229_(_0994_, _0993_, _0794_);
    or _3230_(_0415_, _0994_, _0987_);
    and _3231_(_0995_, _0792_, state[25]);
    xor _3232_(_0996_, round_key[25], state[25]);
    and _3233_(_0997_, _0996_, _0779_);
    and _3234_(_0998_, _0997_, encrypting);
    and _3235_(_0999_, _0998_, _0781_);
    and _3236_(_1000_, _0799_, plaintext[25]);
    or _3237_(_1001_, _1000_, _0999_);
    and _3238_(_1002_, _1001_, _0794_);
    or _3239_(_0416_, _1002_, _0995_);
    and _3240_(_1003_, _0792_, state[26]);
    xor _3241_(_1004_, round_key[26], state[26]);
    and _3242_(_1005_, _1004_, _0779_);
    and _3243_(_1006_, _1005_, encrypting);
    and _3244_(_1007_, _1006_, _0781_);
    and _3245_(_1008_, _0799_, plaintext[26]);
    or _3246_(_1009_, _1008_, _1007_);
    and _3247_(_1010_, _1009_, _0794_);
    or _3248_(_0417_, _1010_, _1003_);
    and _3249_(_1011_, _0792_, state[27]);
    xor _3250_(_1012_, round_key[27], state[27]);
    and _3251_(_1013_, _1012_, _0779_);
    and _3252_(_1014_, _1013_, encrypting);
    and _3253_(_1015_, _1014_, _0781_);
    and _3254_(_1016_, _0799_, plaintext[27]);
    or _3255_(_1017_, _1016_, _1015_);
    and _3256_(_1018_, _1017_, _0794_);
    or _3257_(_0418_, _1018_, _1011_);
    and _3258_(_1019_, _0792_, state[28]);
    xor _3259_(_1020_, round_key[28], state[28]);
    and _3260_(_1021_, _1020_, _0779_);
    and _3261_(_1022_, _1021_, encrypting);
    and _3262_(_1023_, _1022_, _0781_);
    and _3263_(_1024_, _0799_, plaintext[28]);
    or _3264_(_1025_, _1024_, _1023_);
    and _3265_(_1026_, _1025_, _0794_);
    or _3266_(_0419_, _1026_, _1019_);
    and _3267_(_1027_, _0792_, state[29]);
    xor _3268_(_1028_, round_key[29], state[29]);
    and _3269_(_1029_, _1028_, _0779_);
    and _3270_(_1030_, _1029_, encrypting);
    and _3271_(_1031_, _1030_, _0781_);
    and _3272_(_1032_, _0799_, plaintext[29]);
    or _3273_(_1033_, _1032_, _1031_);
    and _3274_(_1034_, _1033_, _0794_);
    or _3275_(_0420_, _1034_, _1027_);
    and _3276_(_1035_, _0792_, state[30]);
    xor _3277_(_1036_, round_key[30], state[30]);
    and _3278_(_1037_, _1036_, _0779_);
    and _3279_(_1038_, _1037_, encrypting);
    and _3280_(_1039_, _1038_, _0781_);
    and _3281_(_1040_, _0799_, plaintext[30]);
    or _3282_(_1041_, _1040_, _1039_);
    and _3283_(_1042_, _1041_, _0794_);
    or _3284_(_0421_, _1042_, _1035_);
    and _3285_(_1043_, _0792_, state[31]);
    xor _3286_(_1044_, round_key[31], state[31]);
    and _3287_(_1045_, _1044_, _0779_);
    and _3288_(_1046_, _1045_, encrypting);
    and _3289_(_1047_, _1046_, _0781_);
    and _3290_(_1048_, _0799_, plaintext[31]);
    or _3291_(_1049_, _1048_, _1047_);
    and _3292_(_1050_, _1049_, _0794_);
    or _3293_(_0422_, _1050_, _1043_);
    and _3294_(_1051_, _0792_, state[32]);
    xor _3295_(_1052_, round_key[32], state[32]);
    and _3296_(_1053_, _1052_, _0779_);
    and _3297_(_1054_, _1053_, encrypting);
    and _3298_(_1055_, _1054_, _0781_);
    and _3299_(_1056_, _0799_, plaintext[32]);
    or _3300_(_1057_, _1056_, _1055_);
    and _3301_(_1058_, _1057_, _0794_);
    or _3302_(_0423_, _1058_, _1051_);
    and _3303_(_1059_, _0792_, state[33]);
    xor _3304_(_1060_, round_key[33], state[33]);
    and _3305_(_1061_, _1060_, _0779_);
    and _3306_(_1062_, _1061_, encrypting);
    and _3307_(_1063_, _1062_, _0781_);
    and _3308_(_1064_, _0799_, plaintext[33]);
    or _3309_(_1065_, _1064_, _1063_);
    and _3310_(_1066_, _1065_, _0794_);
    or _3311_(_0424_, _1066_, _1059_);
    and _3312_(_1067_, _0792_, state[34]);
    xor _3313_(_1068_, round_key[34], state[34]);
    and _3314_(_1069_, _1068_, _0779_);
    and _3315_(_1070_, _1069_, encrypting);
    and _3316_(_1071_, _1070_, _0781_);
    and _3317_(_1072_, _0799_, plaintext[34]);
    or _3318_(_1073_, _1072_, _1071_);
    and _3319_(_1074_, _1073_, _0794_);
    or _3320_(_0425_, _1074_, _1067_);
    and _3321_(_1075_, _0792_, state[35]);
    xor _3322_(_1076_, round_key[35], state[35]);
    and _3323_(_1077_, _1076_, _0779_);
    and _3324_(_1078_, _1077_, encrypting);
    and _3325_(_1079_, _1078_, _0781_);
    and _3326_(_1080_, _0799_, plaintext[35]);
    or _3327_(_1081_, _1080_, _1079_);
    and _3328_(_1082_, _1081_, _0794_);
    or _3329_(_0426_, _1082_, _1075_);
    and _3330_(_1083_, _0792_, state[36]);
    xor _3331_(_1084_, round_key[36], state[36]);
    and _3332_(_1085_, _1084_, _0779_);
    and _3333_(_1086_, _1085_, encrypting);
    and _3334_(_1087_, _1086_, _0781_);
    and _3335_(_1088_, _0799_, plaintext[36]);
    or _3336_(_1089_, _1088_, _1087_);
    and _3337_(_1090_, _1089_, _0794_);
    or _3338_(_0427_, _1090_, _1083_);
    and _3339_(_1091_, _0792_, state[37]);
    xor _3340_(_1092_, round_key[37], state[37]);
    and _3341_(_1093_, _1092_, _0779_);
    and _3342_(_1094_, _1093_, encrypting);
    and _3343_(_1095_, _1094_, _0781_);
    and _3344_(_1096_, _0799_, plaintext[37]);
    or _3345_(_1097_, _1096_, _1095_);
    and _3346_(_1098_, _1097_, _0794_);
    or _3347_(_0428_, _1098_, _1091_);
    and _3348_(_1099_, _0792_, state[38]);
    xor _3349_(_1100_, round_key[38], state[38]);
    and _3350_(_1101_, _1100_, _0779_);
    and _3351_(_1102_, _1101_, encrypting);
    and _3352_(_1103_, _1102_, _0781_);
    and _3353_(_1104_, _0799_, plaintext[38]);
    or _3354_(_1105_, _1104_, _1103_);
    and _3355_(_1106_, _1105_, _0794_);
    or _3356_(_0429_, _1106_, _1099_);
    and _3357_(_1107_, _0792_, state[39]);
    xor _3358_(_1108_, round_key[39], state[39]);
    and _3359_(_1109_, _1108_, _0779_);
    and _3360_(_1110_, _1109_, encrypting);
    and _3361_(_1111_, _1110_, _0781_);
    and _3362_(_1112_, _0799_, plaintext[39]);
    or _3363_(_1113_, _1112_, _1111_);
    and _3364_(_1114_, _1113_, _0794_);
    or _3365_(_0430_, _1114_, _1107_);
    and _3366_(_1115_, _0792_, state[40]);
    xor _3367_(_1116_, round_key[40], state[40]);
    and _3368_(_1117_, _1116_, _0779_);
    and _3369_(_1118_, _1117_, encrypting);
    and _3370_(_1119_, _1118_, _0781_);
    and _3371_(_1120_, _0799_, plaintext[40]);
    or _3372_(_1121_, _1120_, _1119_);
    and _3373_(_1122_, _1121_, _0794_);
    or _3374_(_0431_, _1122_, _1115_);
    and _3375_(_1123_, _0792_, state[41]);
    xor _3376_(_1124_, round_key[41], state[41]);
    and _3377_(_1125_, _1124_, _0779_);
    and _3378_(_1126_, _1125_, encrypting);
    and _3379_(_1127_, _1126_, _0781_);
    and _3380_(_1128_, _0799_, plaintext[41]);
    or _3381_(_1129_, _1128_, _1127_);
    and _3382_(_1130_, _1129_, _0794_);
    or _3383_(_0432_, _1130_, _1123_);
    and _3384_(_1131_, _0792_, state[42]);
    xor _3385_(_1132_, round_key[42], state[42]);
    and _3386_(_1133_, _1132_, _0779_);
    and _3387_(_1134_, _1133_, encrypting);
    and _3388_(_1135_, _1134_, _0781_);
    and _3389_(_1136_, _0799_, plaintext[42]);
    or _3390_(_1137_, _1136_, _1135_);
    and _3391_(_1138_, _1137_, _0794_);
    or _3392_(_0433_, _1138_, _1131_);
    and _3393_(_1139_, _0792_, state[43]);
    xor _3394_(_1140_, round_key[43], state[43]);
    and _3395_(_1141_, _1140_, _0779_);
    and _3396_(_1142_, _1141_, encrypting);
    and _3397_(_1143_, _1142_, _0781_);
    and _3398_(_1144_, _0799_, plaintext[43]);
    or _3399_(_1145_, _1144_, _1143_);
    and _3400_(_1146_, _1145_, _0794_);
    or _3401_(_0434_, _1146_, _1139_);
    and _3402_(_1147_, _0792_, state[44]);
    xor _3403_(_1148_, round_key[44], state[44]);
    and _3404_(_1149_, _1148_, _0779_);
    and _3405_(_1150_, _1149_, encrypting);
    and _3406_(_1151_, _1150_, _0781_);
    and _3407_(_1152_, _0799_, plaintext[44]);
    or _3408_(_1153_, _1152_, _1151_);
    and _3409_(_1154_, _1153_, _0794_);
    or _3410_(_0435_, _1154_, _1147_);
    and _3411_(_1155_, _0792_, state[45]);
    xor _3412_(_1156_, round_key[45], state[45]);
    and _3413_(_1157_, _1156_, _0779_);
    and _3414_(_1158_, _1157_, encrypting);
    and _3415_(_1159_, _1158_, _0781_);
    and _3416_(_1160_, _0799_, plaintext[45]);
    or _3417_(_1161_, _1160_, _1159_);
    and _3418_(_1162_, _1161_, _0794_);
    or _3419_(_0436_, _1162_, _1155_);
    and _3420_(_1163_, _0792_, state[46]);
    xor _3421_(_1164_, round_key[46], state[46]);
    and _3422_(_1165_, _1164_, _0779_);
    and _3423_(_1166_, _1165_, encrypting);
    and _3424_(_1167_, _1166_, _0781_);
    and _3425_(_1168_, _0799_, plaintext[46]);
    or _3426_(_1169_, _1168_, _1167_);
    and _3427_(_1170_, _1169_, _0794_);
    or _3428_(_0437_, _1170_, _1163_);
    and _3429_(_1171_, _0792_, state[47]);
    xor _3430_(_1172_, round_key[47], state[47]);
    and _3431_(_1173_, _1172_, _0779_);
    and _3432_(_1174_, _1173_, encrypting);
    and _3433_(_1175_, _1174_, _0781_);
    and _3434_(_1176_, _0799_, plaintext[47]);
    or _3435_(_1177_, _1176_, _1175_);
    and _3436_(_1178_, _1177_, _0794_);
    or _3437_(_0438_, _1178_, _1171_);
    and _3438_(_1179_, _0792_, state[48]);
    xor _3439_(_1180_, round_key[48], state[48]);
    and _3440_(_1181_, _1180_, _0779_);
    and _3441_(_1182_, _1181_, encrypting);
    and _3442_(_1183_, _1182_, _0781_);
    and _3443_(_1184_, _0799_, plaintext[48]);
    or _3444_(_1185_, _1184_, _1183_);
    and _3445_(_1186_, _1185_, _0794_);
    or _3446_(_0439_, _1186_, _1179_);
    and _3447_(_1187_, _0792_, state[49]);
    xor _3448_(_1188_, round_key[49], state[49]);
    and _3449_(_1189_, _1188_, _0779_);
    and _3450_(_1190_, _1189_, encrypting);
    and _3451_(_1191_, _1190_, _0781_);
    and _3452_(_1192_, _0799_, plaintext[49]);
    or _3453_(_1193_, _1192_, _1191_);
    and _3454_(_1194_, _1193_, _0794_);
    or _3455_(_0440_, _1194_, _1187_);
    and _3456_(_1195_, _0792_, state[50]);
    xor _3457_(_1196_, round_key[50], state[50]);
    and _3458_(_1197_, _1196_, _0779_);
    and _3459_(_1198_, _1197_, encrypting);
    and _3460_(_1199_, _1198_, _0781_);
    and _3461_(_1200_, _0799_, plaintext[50]);
    or _3462_(_1201_, _1200_, _1199_);
    and _3463_(_1202_, _1201_, _0794_);
    or _3464_(_0441_, _1202_, _1195_);
    and _3465_(_1203_, _0792_, state[51]);
    xor _3466_(_1204_, round_key[51], state[51]);
    and _3467_(_1205_, _1204_, _0779_);
    and _3468_(_1206_, _1205_, encrypting);
    and _3469_(_1207_, _1206_, _0781_);
    and _3470_(_1208_, _0799_, plaintext[51]);
    or _3471_(_1209_, _1208_, _1207_);
    and _3472_(_1210_, _1209_, _0794_);
    or _3473_(_0442_, _1210_, _1203_);
    and _3474_(_1211_, _0792_, state[52]);
    xor _3475_(_1212_, round_key[52], state[52]);
    and _3476_(_1213_, _1212_, _0779_);
    and _3477_(_1214_, _1213_, encrypting);
    and _3478_(_1215_, _1214_, _0781_);
    and _3479_(_1216_, _0799_, plaintext[52]);
    or _3480_(_1217_, _1216_, _1215_);
    and _3481_(_1218_, _1217_, _0794_);
    or _3482_(_0443_, _1218_, _1211_);
    and _3483_(_1219_, _0792_, state[53]);
    xor _3484_(_1220_, round_key[53], state[53]);
    and _3485_(_1221_, _1220_, _0779_);
    and _3486_(_1222_, _1221_, encrypting);
    and _3487_(_1223_, _1222_, _0781_);
    and _3488_(_1224_, _0799_, plaintext[53]);
    or _3489_(_1225_, _1224_, _1223_);
    and _3490_(_1226_, _1225_, _0794_);
    or _3491_(_0444_, _1226_, _1219_);
    and _3492_(_1227_, _0792_, state[54]);
    xor _3493_(_1228_, round_key[54], state[54]);
    and _3494_(_1229_, _1228_, _0779_);
    and _3495_(_1230_, _1229_, encrypting);
    and _3496_(_1231_, _1230_, _0781_);
    and _3497_(_1232_, _0799_, plaintext[54]);
    or _3498_(_1233_, _1232_, _1231_);
    and _3499_(_1234_, _1233_, _0794_);
    or _3500_(_0445_, _1234_, _1227_);
    and _3501_(_1235_, _0792_, state[55]);
    xor _3502_(_1236_, round_key[55], state[55]);
    and _3503_(_1237_, _1236_, _0779_);
    and _3504_(_1238_, _1237_, encrypting);
    and _3505_(_1239_, _1238_, _0781_);
    and _3506_(_1240_, _0799_, plaintext[55]);
    or _3507_(_1241_, _1240_, _1239_);
    and _3508_(_1242_, _1241_, _0794_);
    or _3509_(_0446_, _1242_, _1235_);
    and _3510_(_1243_, _0792_, state[56]);
    xor _3511_(_1244_, round_key[56], state[56]);
    and _3512_(_1245_, _1244_, _0779_);
    and _3513_(_1246_, _1245_, encrypting);
    and _3514_(_1247_, _1246_, _0781_);
    and _3515_(_1248_, _0799_, plaintext[56]);
    or _3516_(_1249_, _1248_, _1247_);
    and _3517_(_1250_, _1249_, _0794_);
    or _3518_(_0447_, _1250_, _1243_);
    and _3519_(_1251_, _0792_, state[57]);
    xor _3520_(_1252_, round_key[57], state[57]);
    and _3521_(_1253_, _1252_, _0779_);
    and _3522_(_1254_, _1253_, encrypting);
    and _3523_(_1255_, _1254_, _0781_);
    and _3524_(_1256_, _0799_, plaintext[57]);
    or _3525_(_1257_, _1256_, _1255_);
    and _3526_(_1258_, _1257_, _0794_);
    or _3527_(_0448_, _1258_, _1251_);
    and _3528_(_1259_, _0792_, state[58]);
    xor _3529_(_1260_, round_key[58], state[58]);
    and _3530_(_1261_, _1260_, _0779_);
    and _3531_(_1262_, _1261_, encrypting);
    and _3532_(_1263_, _1262_, _0781_);
    and _3533_(_1264_, _0799_, plaintext[58]);
    or _3534_(_1265_, _1264_, _1263_);
    and _3535_(_1266_, _1265_, _0794_);
    or _3536_(_0449_, _1266_, _1259_);
    and _3537_(_1267_, _0792_, state[59]);
    xor _3538_(_1268_, round_key[59], state[59]);
    and _3539_(_1269_, _1268_, _0779_);
    and _3540_(_1270_, _1269_, encrypting);
    and _3541_(_1271_, _1270_, _0781_);
    and _3542_(_1272_, _0799_, plaintext[59]);
    or _3543_(_1273_, _1272_, _1271_);
    and _3544_(_1274_, _1273_, _0794_);
    or _3545_(_0450_, _1274_, _1267_);
    and _3546_(_1275_, _0792_, state[60]);
    xor _3547_(_1276_, round_key[60], state[60]);
    and _3548_(_1277_, _1276_, _0779_);
    and _3549_(_1278_, _1277_, encrypting);
    and _3550_(_1279_, _1278_, _0781_);
    and _3551_(_1280_, _0799_, plaintext[60]);
    or _3552_(_1281_, _1280_, _1279_);
    and _3553_(_1282_, _1281_, _0794_);
    or _3554_(_0451_, _1282_, _1275_);
    and _3555_(_1283_, _0792_, state[61]);
    xor _3556_(_1284_, round_key[61], state[61]);
    and _3557_(_1285_, _1284_, _0779_);
    and _3558_(_1286_, _1285_, encrypting);
    and _3559_(_1287_, _1286_, _0781_);
    and _3560_(_1288_, _0799_, plaintext[61]);
    or _3561_(_1289_, _1288_, _1287_);
    and _3562_(_1290_, _1289_, _0794_);
    or _3563_(_0452_, _1290_, _1283_);
    and _3564_(_1291_, _0792_, state[62]);
    xor _3565_(_1292_, round_key[62], state[62]);
    and _3566_(_1293_, _1292_, _0779_);
    and _3567_(_1294_, _1293_, encrypting);
    and _3568_(_1295_, _1294_, _0781_);
    and _3569_(_1296_, _0799_, plaintext[62]);
    or _3570_(_1297_, _1296_, _1295_);
    and _3571_(_1298_, _1297_, _0794_);
    or _3572_(_0453_, _1298_, _1291_);
    and _3573_(_1299_, _0792_, state[63]);
    xor _3574_(_1300_, round_key[63], state[63]);
    and _3575_(_1301_, _1300_, _0779_);
    and _3576_(_1302_, _1301_, encrypting);
    and _3577_(_1303_, _1302_, _0781_);
    and _3578_(_1304_, _0799_, plaintext[63]);
    or _3579_(_1305_, _1304_, _1303_);
    and _3580_(_1306_, _1305_, _0794_);
    or _3581_(_0454_, _1306_, _1299_);
    and _3582_(_1307_, _0792_, state[64]);
    xor _3583_(_1308_, round_key[64], state[64]);
    and _3584_(_1309_, _1308_, _0779_);
    and _3585_(_1310_, _1309_, encrypting);
    and _3586_(_1311_, _1310_, _0781_);
    and _3587_(_1312_, _0799_, plaintext[64]);
    or _3588_(_1313_, _1312_, _1311_);
    and _3589_(_1314_, _1313_, _0794_);
    or _3590_(_0455_, _1314_, _1307_);
    and _3591_(_1315_, _0792_, state[65]);
    xor _3592_(_1316_, round_key[65], state[65]);
    and _3593_(_1317_, _1316_, _0779_);
    and _3594_(_1318_, _1317_, encrypting);
    and _3595_(_1319_, _1318_, _0781_);
    and _3596_(_1320_, _0799_, plaintext[65]);
    or _3597_(_1321_, _1320_, _1319_);
    and _3598_(_1322_, _1321_, _0794_);
    or _3599_(_0456_, _1322_, _1315_);
    and _3600_(_1323_, _0792_, state[66]);
    xor _3601_(_1324_, round_key[66], state[66]);
    and _3602_(_1325_, _1324_, _0779_);
    and _3603_(_1326_, _1325_, encrypting);
    and _3604_(_1327_, _1326_, _0781_);
    and _3605_(_1328_, _0799_, plaintext[66]);
    or _3606_(_1329_, _1328_, _1327_);
    and _3607_(_1330_, _1329_, _0794_);
    or _3608_(_0457_, _1330_, _1323_);
    and _3609_(_1331_, _0792_, state[67]);
    xor _3610_(_1332_, round_key[67], state[67]);
    and _3611_(_1333_, _1332_, _0779_);
    and _3612_(_1334_, _1333_, encrypting);
    and _3613_(_1335_, _1334_, _0781_);
    and _3614_(_1336_, _0799_, plaintext[67]);
    or _3615_(_1337_, _1336_, _1335_);
    and _3616_(_1338_, _1337_, _0794_);
    or _3617_(_0458_, _1338_, _1331_);
    and _3618_(_1339_, _0792_, state[68]);
    xor _3619_(_1340_, round_key[68], state[68]);
    and _3620_(_1341_, _1340_, _0779_);
    and _3621_(_1342_, _1341_, encrypting);
    and _3622_(_1343_, _1342_, _0781_);
    and _3623_(_1344_, _0799_, plaintext[68]);
    or _3624_(_1345_, _1344_, _1343_);
    and _3625_(_1346_, _1345_, _0794_);
    or _3626_(_0459_, _1346_, _1339_);
    and _3627_(_1347_, _0792_, state[69]);
    xor _3628_(_1348_, round_key[69], state[69]);
    and _3629_(_1349_, _1348_, _0779_);
    and _3630_(_1350_, _1349_, encrypting);
    and _3631_(_1351_, _1350_, _0781_);
    and _3632_(_1352_, _0799_, plaintext[69]);
    or _3633_(_1353_, _1352_, _1351_);
    and _3634_(_1354_, _1353_, _0794_);
    or _3635_(_0460_, _1354_, _1347_);
    and _3636_(_1355_, _0792_, state[70]);
    xor _3637_(_1356_, round_key[70], state[70]);
    and _3638_(_1357_, _1356_, _0779_);
    and _3639_(_1358_, _1357_, encrypting);
    and _3640_(_1359_, _1358_, _0781_);
    and _3641_(_1360_, _0799_, plaintext[70]);
    or _3642_(_1361_, _1360_, _1359_);
    and _3643_(_1362_, _1361_, _0794_);
    or _3644_(_0461_, _1362_, _1355_);
    and _3645_(_1363_, _0792_, state[71]);
    xor _3646_(_1364_, round_key[71], state[71]);
    and _3647_(_1365_, _1364_, _0779_);
    and _3648_(_1366_, _1365_, encrypting);
    and _3649_(_1367_, _1366_, _0781_);
    and _3650_(_1368_, _0799_, plaintext[71]);
    or _3651_(_1369_, _1368_, _1367_);
    and _3652_(_1370_, _1369_, _0794_);
    or _3653_(_0462_, _1370_, _1363_);
    and _3654_(_1371_, _0792_, state[72]);
    xor _3655_(_1372_, round_key[72], state[72]);
    and _3656_(_1373_, _1372_, _0779_);
    and _3657_(_1374_, _1373_, encrypting);
    and _3658_(_1375_, _1374_, _0781_);
    and _3659_(_1376_, _0799_, plaintext[72]);
    or _3660_(_1377_, _1376_, _1375_);
    and _3661_(_1378_, _1377_, _0794_);
    or _3662_(_0463_, _1378_, _1371_);
    and _3663_(_1379_, _0792_, state[73]);
    xor _3664_(_1380_, round_key[73], state[73]);
    and _3665_(_1381_, _1380_, _0779_);
    and _3666_(_1382_, _1381_, encrypting);
    and _3667_(_1383_, _1382_, _0781_);
    and _3668_(_1384_, _0799_, plaintext[73]);
    or _3669_(_1385_, _1384_, _1383_);
    and _3670_(_1386_, _1385_, _0794_);
    or _3671_(_0464_, _1386_, _1379_);
    and _3672_(_1387_, _0792_, state[74]);
    xor _3673_(_1388_, round_key[74], state[74]);
    and _3674_(_1389_, _1388_, _0779_);
    and _3675_(_1390_, _1389_, encrypting);
    and _3676_(_1391_, _1390_, _0781_);
    and _3677_(_1392_, _0799_, plaintext[74]);
    or _3678_(_1393_, _1392_, _1391_);
    and _3679_(_1394_, _1393_, _0794_);
    or _3680_(_0465_, _1394_, _1387_);
    and _3681_(_1395_, _0792_, state[75]);
    xor _3682_(_1396_, round_key[75], state[75]);
    and _3683_(_1397_, _1396_, _0779_);
    and _3684_(_1398_, _1397_, encrypting);
    and _3685_(_1399_, _1398_, _0781_);
    and _3686_(_1400_, _0799_, plaintext[75]);
    or _3687_(_1401_, _1400_, _1399_);
    and _3688_(_1402_, _1401_, _0794_);
    or _3689_(_0466_, _1402_, _1395_);
    and _3690_(_1403_, _0792_, state[76]);
    xor _3691_(_1404_, round_key[76], state[76]);
    and _3692_(_1405_, _1404_, _0779_);
    and _3693_(_1406_, _1405_, encrypting);
    and _3694_(_1407_, _1406_, _0781_);
    and _3695_(_1408_, _0799_, plaintext[76]);
    or _3696_(_1409_, _1408_, _1407_);
    and _3697_(_1410_, _1409_, _0794_);
    or _3698_(_0467_, _1410_, _1403_);
    and _3699_(_1411_, _0792_, state[77]);
    xor _3700_(_1412_, round_key[77], state[77]);
    and _3701_(_1413_, _1412_, _0779_);
    and _3702_(_1414_, _1413_, encrypting);
    and _3703_(_1415_, _1414_, _0781_);
    and _3704_(_1416_, _0799_, plaintext[77]);
    or _3705_(_1417_, _1416_, _1415_);
    and _3706_(_1418_, _1417_, _0794_);
    or _3707_(_0468_, _1418_, _1411_);
    and _3708_(_1419_, _0792_, state[78]);
    xor _3709_(_1420_, round_key[78], state[78]);
    and _3710_(_1421_, _1420_, _0779_);
    and _3711_(_1422_, _1421_, encrypting);
    and _3712_(_1423_, _1422_, _0781_);
    and _3713_(_1424_, _0799_, plaintext[78]);
    or _3714_(_1425_, _1424_, _1423_);
    and _3715_(_1426_, _1425_, _0794_);
    or _3716_(_0469_, _1426_, _1419_);
    and _3717_(_1427_, _0792_, state[79]);
    xor _3718_(_1428_, round_key[79], state[79]);
    and _3719_(_1429_, _1428_, _0779_);
    and _3720_(_1430_, _1429_, encrypting);
    and _3721_(_1431_, _1430_, _0781_);
    and _3722_(_1432_, _0799_, plaintext[79]);
    or _3723_(_1433_, _1432_, _1431_);
    and _3724_(_1434_, _1433_, _0794_);
    or _3725_(_0470_, _1434_, _1427_);
    and _3726_(_1435_, _0792_, state[80]);
    xor _3727_(_1436_, round_key[80], state[80]);
    and _3728_(_1437_, _1436_, _0779_);
    and _3729_(_1438_, _1437_, encrypting);
    and _3730_(_1439_, _1438_, _0781_);
    and _3731_(_1440_, _0799_, plaintext[80]);
    or _3732_(_1441_, _1440_, _1439_);
    and _3733_(_1442_, _1441_, _0794_);
    or _3734_(_0471_, _1442_, _1435_);
    and _3735_(_1443_, _0792_, state[81]);
    xor _3736_(_1444_, round_key[81], state[81]);
    and _3737_(_1445_, _1444_, _0779_);
    and _3738_(_1446_, _1445_, encrypting);
    and _3739_(_1447_, _1446_, _0781_);
    and _3740_(_1448_, _0799_, plaintext[81]);
    or _3741_(_1449_, _1448_, _1447_);
    and _3742_(_1450_, _1449_, _0794_);
    or _3743_(_0472_, _1450_, _1443_);
    and _3744_(_1451_, _0792_, state[82]);
    xor _3745_(_1452_, round_key[82], state[82]);
    and _3746_(_1453_, _1452_, _0779_);
    and _3747_(_1454_, _1453_, encrypting);
    and _3748_(_1455_, _1454_, _0781_);
    and _3749_(_1456_, _0799_, plaintext[82]);
    or _3750_(_1457_, _1456_, _1455_);
    and _3751_(_1458_, _1457_, _0794_);
    or _3752_(_0473_, _1458_, _1451_);
    and _3753_(_1459_, _0792_, state[83]);
    xor _3754_(_1460_, round_key[83], state[83]);
    and _3755_(_1461_, _1460_, _0779_);
    and _3756_(_1462_, _1461_, encrypting);
    and _3757_(_1463_, _1462_, _0781_);
    and _3758_(_1464_, _0799_, plaintext[83]);
    or _3759_(_1465_, _1464_, _1463_);
    and _3760_(_1466_, _1465_, _0794_);
    or _3761_(_0474_, _1466_, _1459_);
    and _3762_(_1467_, _0792_, state[84]);
    xor _3763_(_1468_, round_key[84], state[84]);
    and _3764_(_1469_, _1468_, _0779_);
    and _3765_(_1470_, _1469_, encrypting);
    and _3766_(_1471_, _1470_, _0781_);
    and _3767_(_1472_, _0799_, plaintext[84]);
    or _3768_(_1473_, _1472_, _1471_);
    and _3769_(_1474_, _1473_, _0794_);
    or _3770_(_0475_, _1474_, _1467_);
    and _3771_(_1475_, _0792_, state[85]);
    xor _3772_(_1476_, round_key[85], state[85]);
    and _3773_(_1477_, _1476_, _0779_);
    and _3774_(_1478_, _1477_, encrypting);
    and _3775_(_1479_, _1478_, _0781_);
    and _3776_(_1480_, _0799_, plaintext[85]);
    or _3777_(_1481_, _1480_, _1479_);
    and _3778_(_1482_, _1481_, _0794_);
    or _3779_(_0476_, _1482_, _1475_);
    and _3780_(_1483_, _0792_, state[86]);
    xor _3781_(_1484_, round_key[86], state[86]);
    and _3782_(_1485_, _1484_, _0779_);
    and _3783_(_1486_, _1485_, encrypting);
    and _3784_(_1487_, _1486_, _0781_);
    and _3785_(_1488_, _0799_, plaintext[86]);
    or _3786_(_1489_, _1488_, _1487_);
    and _3787_(_1490_, _1489_, _0794_);
    or _3788_(_0477_, _1490_, _1483_);
    and _3789_(_1491_, _0792_, state[87]);
    xor _3790_(_1492_, round_key[87], state[87]);
    and _3791_(_1493_, _1492_, _0779_);
    and _3792_(_1494_, _1493_, encrypting);
    and _3793_(_1495_, _1494_, _0781_);
    and _3794_(_1496_, _0799_, plaintext[87]);
    or _3795_(_1497_, _1496_, _1495_);
    and _3796_(_1498_, _1497_, _0794_);
    or _3797_(_0478_, _1498_, _1491_);
    and _3798_(_1499_, _0792_, state[88]);
    xor _3799_(_1500_, round_key[88], state[88]);
    and _3800_(_1501_, _1500_, _0779_);
    and _3801_(_1502_, _1501_, encrypting);
    and _3802_(_1503_, _1502_, _0781_);
    and _3803_(_1504_, _0799_, plaintext[88]);
    or _3804_(_1505_, _1504_, _1503_);
    and _3805_(_1506_, _1505_, _0794_);
    or _3806_(_0479_, _1506_, _1499_);
    and _3807_(_1507_, _0792_, state[89]);
    xor _3808_(_1508_, round_key[89], state[89]);
    and _3809_(_1509_, _1508_, _0779_);
    and _3810_(_1510_, _1509_, encrypting);
    and _3811_(_1511_, _1510_, _0781_);
    and _3812_(_1512_, _0799_, plaintext[89]);
    or _3813_(_1513_, _1512_, _1511_);
    and _3814_(_1514_, _1513_, _0794_);
    or _3815_(_0480_, _1514_, _1507_);
    and _3816_(_1515_, _0792_, state[90]);
    xor _3817_(_1516_, round_key[90], state[90]);
    and _3818_(_1517_, _1516_, _0779_);
    and _3819_(_1518_, _1517_, encrypting);
    and _3820_(_1519_, _1518_, _0781_);
    and _3821_(_1520_, _0799_, plaintext[90]);
    or _3822_(_1521_, _1520_, _1519_);
    and _3823_(_1522_, _1521_, _0794_);
    or _3824_(_0481_, _1522_, _1515_);
    and _3825_(_1523_, _0792_, state[91]);
    xor _3826_(_1524_, round_key[91], state[91]);
    and _3827_(_1525_, _1524_, _0779_);
    and _3828_(_1526_, _1525_, encrypting);
    and _3829_(_1527_, _1526_, _0781_);
    and _3830_(_1528_, _0799_, plaintext[91]);
    or _3831_(_1529_, _1528_, _1527_);
    and _3832_(_1530_, _1529_, _0794_);
    or _3833_(_0482_, _1530_, _1523_);
    and _3834_(_1531_, _0792_, state[92]);
    xor _3835_(_1532_, round_key[92], state[92]);
    and _3836_(_1533_, _1532_, _0779_);
    and _3837_(_1534_, _1533_, encrypting);
    and _3838_(_1535_, _1534_, _0781_);
    and _3839_(_1536_, _0799_, plaintext[92]);
    or _3840_(_1537_, _1536_, _1535_);
    and _3841_(_1538_, _1537_, _0794_);
    or _3842_(_0483_, _1538_, _1531_);
    and _3843_(_1539_, _0792_, state[93]);
    xor _3844_(_1540_, round_key[93], state[93]);
    and _3845_(_1541_, _1540_, _0779_);
    and _3846_(_1542_, _1541_, encrypting);
    and _3847_(_1543_, _1542_, _0781_);
    and _3848_(_1544_, _0799_, plaintext[93]);
    or _3849_(_1545_, _1544_, _1543_);
    and _3850_(_1546_, _1545_, _0794_);
    or _3851_(_0484_, _1546_, _1539_);
    and _3852_(_1547_, _0792_, state[94]);
    xor _3853_(_1548_, round_key[94], state[94]);
    and _3854_(_1549_, _1548_, _0779_);
    and _3855_(_1550_, _1549_, encrypting);
    and _3856_(_1551_, _1550_, _0781_);
    and _3857_(_1552_, _0799_, plaintext[94]);
    or _3858_(_1553_, _1552_, _1551_);
    and _3859_(_1554_, _1553_, _0794_);
    or _3860_(_0485_, _1554_, _1547_);
    and _3861_(_1555_, _0792_, state[95]);
    xor _3862_(_1556_, round_key[95], state[95]);
    and _3863_(_1557_, _1556_, _0779_);
    and _3864_(_1558_, _1557_, encrypting);
    and _3865_(_1559_, _1558_, _0781_);
    and _3866_(_1560_, _0799_, plaintext[95]);
    or _3867_(_1561_, _1560_, _1559_);
    and _3868_(_1562_, _1561_, _0794_);
    or _3869_(_0486_, _1562_, _1555_);
    and _3870_(_1563_, _0792_, state[96]);
    xor _3871_(_1564_, round_key[96], state[96]);
    and _3872_(_1565_, _1564_, _0779_);
    and _3873_(_1566_, _1565_, encrypting);
    and _3874_(_1567_, _1566_, _0781_);
    and _3875_(_1568_, _0799_, plaintext[96]);
    or _3876_(_1569_, _1568_, _1567_);
    and _3877_(_1570_, _1569_, _0794_);
    or _3878_(_0487_, _1570_, _1563_);
    and _3879_(_1571_, _0792_, state[97]);
    xor _3880_(_1572_, round_key[97], state[97]);
    and _3881_(_1573_, _1572_, _0779_);
    and _3882_(_1574_, _1573_, encrypting);
    and _3883_(_1575_, _1574_, _0781_);
    and _3884_(_1576_, _0799_, plaintext[97]);
    or _3885_(_1577_, _1576_, _1575_);
    and _3886_(_1578_, _1577_, _0794_);
    or _3887_(_0488_, _1578_, _1571_);
    and _3888_(_1579_, _0792_, state[98]);
    xor _3889_(_1580_, round_key[98], state[98]);
    and _3890_(_1581_, _1580_, _0779_);
    and _3891_(_1582_, _1581_, encrypting);
    and _3892_(_1583_, _1582_, _0781_);
    and _3893_(_1584_, _0799_, plaintext[98]);
    or _3894_(_1585_, _1584_, _1583_);
    and _3895_(_1586_, _1585_, _0794_);
    or _3896_(_0489_, _1586_, _1579_);
    and _3897_(_1587_, _0792_, state[99]);
    xor _3898_(_1588_, round_key[99], state[99]);
    and _3899_(_1589_, _1588_, _0779_);
    and _3900_(_1590_, _1589_, encrypting);
    and _3901_(_1591_, _1590_, _0781_);
    and _3902_(_1592_, _0799_, plaintext[99]);
    or _3903_(_1593_, _1592_, _1591_);
    and _3904_(_1594_, _1593_, _0794_);
    or _3905_(_0490_, _1594_, _1587_);
    and _3906_(_1595_, _0792_, state[100]);
    xor _3907_(_1596_, round_key[100], state[100]);
    and _3908_(_1597_, _1596_, _0779_);
    and _3909_(_1598_, _1597_, encrypting);
    and _3910_(_1599_, _1598_, _0781_);
    and _3911_(_1600_, _0799_, plaintext[100]);
    or _3912_(_1601_, _1600_, _1599_);
    and _3913_(_1602_, _1601_, _0794_);
    or _3914_(_0491_, _1602_, _1595_);
    and _3915_(_1603_, _0792_, state[101]);
    xor _3916_(_1604_, round_key[101], state[101]);
    and _3917_(_1605_, _1604_, _0779_);
    and _3918_(_1606_, _1605_, encrypting);
    and _3919_(_1607_, _1606_, _0781_);
    and _3920_(_1608_, _0799_, plaintext[101]);
    or _3921_(_1609_, _1608_, _1607_);
    and _3922_(_1610_, _1609_, _0794_);
    or _3923_(_0492_, _1610_, _1603_);
    and _3924_(_1611_, _0792_, state[102]);
    xor _3925_(_1612_, round_key[102], state[102]);
    and _3926_(_1613_, _1612_, _0779_);
    and _3927_(_1614_, _1613_, encrypting);
    and _3928_(_1615_, _1614_, _0781_);
    and _3929_(_1616_, _0799_, plaintext[102]);
    or _3930_(_1617_, _1616_, _1615_);
    and _3931_(_1618_, _1617_, _0794_);
    or _3932_(_0493_, _1618_, _1611_);
    and _3933_(_1619_, _0792_, state[103]);
    xor _3934_(_1620_, round_key[103], state[103]);
    and _3935_(_1621_, _1620_, _0779_);
    and _3936_(_1622_, _1621_, encrypting);
    and _3937_(_1623_, _1622_, _0781_);
    and _3938_(_1624_, _0799_, plaintext[103]);
    or _3939_(_1625_, _1624_, _1623_);
    and _3940_(_1626_, _1625_, _0794_);
    or _3941_(_0494_, _1626_, _1619_);
    and _3942_(_1627_, _0792_, state[104]);
    xor _3943_(_1628_, round_key[104], state[104]);
    and _3944_(_1629_, _1628_, _0779_);
    and _3945_(_1630_, _1629_, encrypting);
    and _3946_(_1631_, _1630_, _0781_);
    and _3947_(_1632_, _0799_, plaintext[104]);
    or _3948_(_1633_, _1632_, _1631_);
    and _3949_(_1634_, _1633_, _0794_);
    or _3950_(_0495_, _1634_, _1627_);
    and _3951_(_1635_, _0792_, state[105]);
    xor _3952_(_1636_, round_key[105], state[105]);
    and _3953_(_1637_, _1636_, _0779_);
    and _3954_(_1638_, _1637_, encrypting);
    and _3955_(_1639_, _1638_, _0781_);
    and _3956_(_1640_, _0799_, plaintext[105]);
    or _3957_(_1641_, _1640_, _1639_);
    and _3958_(_1642_, _1641_, _0794_);
    or _3959_(_0496_, _1642_, _1635_);
    and _3960_(_1643_, _0792_, state[106]);
    xor _3961_(_1644_, round_key[106], state[106]);
    and _3962_(_1645_, _1644_, _0779_);
    and _3963_(_1646_, _1645_, encrypting);
    and _3964_(_1647_, _1646_, _0781_);
    and _3965_(_1648_, _0799_, plaintext[106]);
    or _3966_(_1649_, _1648_, _1647_);
    and _3967_(_1650_, _1649_, _0794_);
    or _3968_(_0497_, _1650_, _1643_);
    and _3969_(_1651_, _0792_, state[107]);
    xor _3970_(_1652_, round_key[107], state[107]);
    and _3971_(_1653_, _1652_, _0779_);
    and _3972_(_1654_, _1653_, encrypting);
    and _3973_(_1655_, _1654_, _0781_);
    and _3974_(_1656_, _0799_, plaintext[107]);
    or _3975_(_1657_, _1656_, _1655_);
    and _3976_(_1658_, _1657_, _0794_);
    or _3977_(_0498_, _1658_, _1651_);
    and _3978_(_1659_, _0792_, state[108]);
    xor _3979_(_1660_, round_key[108], state[108]);
    and _3980_(_1661_, _1660_, _0779_);
    and _3981_(_1662_, _1661_, encrypting);
    and _3982_(_1663_, _1662_, _0781_);
    and _3983_(_1664_, _0799_, plaintext[108]);
    or _3984_(_1665_, _1664_, _1663_);
    and _3985_(_1666_, _1665_, _0794_);
    or _3986_(_0499_, _1666_, _1659_);
    and _3987_(_1667_, _0792_, state[109]);
    xor _3988_(_1668_, round_key[109], state[109]);
    and _3989_(_1669_, _1668_, _0779_);
    and _3990_(_1670_, _1669_, encrypting);
    and _3991_(_1671_, _1670_, _0781_);
    and _3992_(_1672_, _0799_, plaintext[109]);
    or _3993_(_1673_, _1672_, _1671_);
    and _3994_(_1674_, _1673_, _0794_);
    or _3995_(_0500_, _1674_, _1667_);
    and _3996_(_1675_, _0792_, state[110]);
    xor _3997_(_1676_, round_key[110], state[110]);
    and _3998_(_1677_, _1676_, _0779_);
    and _3999_(_1678_, _1677_, encrypting);
    and _4000_(_1679_, _1678_, _0781_);
    and _4001_(_1680_, _0799_, plaintext[110]);
    or _4002_(_1681_, _1680_, _1679_);
    and _4003_(_1682_, _1681_, _0794_);
    or _4004_(_0501_, _1682_, _1675_);
    and _4005_(_1683_, _0792_, state[111]);
    xor _4006_(_1684_, round_key[111], state[111]);
    and _4007_(_1685_, _1684_, _0779_);
    and _4008_(_1686_, _1685_, encrypting);
    and _4009_(_1687_, _1686_, _0781_);
    and _4010_(_1688_, _0799_, plaintext[111]);
    or _4011_(_1689_, _1688_, _1687_);
    and _4012_(_1690_, _1689_, _0794_);
    or _4013_(_0502_, _1690_, _1683_);
    and _4014_(_1691_, _0792_, state[112]);
    xor _4015_(_1692_, round_key[112], state[112]);
    and _4016_(_1693_, _1692_, _0779_);
    and _4017_(_1694_, _1693_, encrypting);
    and _4018_(_1695_, _1694_, _0781_);
    and _4019_(_1696_, _0799_, plaintext[112]);
    or _4020_(_1697_, _1696_, _1695_);
    and _4021_(_1698_, _1697_, _0794_);
    or _4022_(_0503_, _1698_, _1691_);
    and _4023_(_1699_, _0792_, state[113]);
    xor _4024_(_1700_, round_key[113], state[113]);
    and _4025_(_1701_, _1700_, _0779_);
    and _4026_(_1702_, _1701_, encrypting);
    and _4027_(_1703_, _1702_, _0781_);
    and _4028_(_1704_, _0799_, plaintext[113]);
    or _4029_(_1705_, _1704_, _1703_);
    and _4030_(_1706_, _1705_, _0794_);
    or _4031_(_0504_, _1706_, _1699_);
    and _4032_(_1707_, _0792_, state[114]);
    xor _4033_(_1708_, round_key[114], state[114]);
    and _4034_(_1709_, _1708_, _0779_);
    and _4035_(_1710_, _1709_, encrypting);
    and _4036_(_1711_, _1710_, _0781_);
    and _4037_(_1712_, _0799_, plaintext[114]);
    or _4038_(_1713_, _1712_, _1711_);
    and _4039_(_1714_, _1713_, _0794_);
    or _4040_(_0505_, _1714_, _1707_);
    and _4041_(_1715_, _0792_, state[115]);
    xor _4042_(_1716_, round_key[115], state[115]);
    and _4043_(_1717_, _1716_, _0779_);
    and _4044_(_1718_, _1717_, encrypting);
    and _4045_(_1719_, _1718_, _0781_);
    and _4046_(_1720_, _0799_, plaintext[115]);
    or _4047_(_1721_, _1720_, _1719_);
    and _4048_(_1722_, _1721_, _0794_);
    or _4049_(_0506_, _1722_, _1715_);
    and _4050_(_1723_, _0792_, state[116]);
    xor _4051_(_1724_, round_key[116], state[116]);
    and _4052_(_1725_, _1724_, _0779_);
    and _4053_(_1726_, _1725_, encrypting);
    and _4054_(_1727_, _1726_, _0781_);
    and _4055_(_1728_, _0799_, plaintext[116]);
    or _4056_(_1729_, _1728_, _1727_);
    and _4057_(_1730_, _1729_, _0794_);
    or _4058_(_0507_, _1730_, _1723_);
    and _4059_(_1731_, _0792_, state[117]);
    xor _4060_(_1732_, round_key[117], state[117]);
    and _4061_(_1733_, _1732_, _0779_);
    and _4062_(_1734_, _1733_, encrypting);
    and _4063_(_1735_, _1734_, _0781_);
    and _4064_(_1736_, _0799_, plaintext[117]);
    or _4065_(_1737_, _1736_, _1735_);
    and _4066_(_1738_, _1737_, _0794_);
    or _4067_(_0508_, _1738_, _1731_);
    and _4068_(_1739_, _0792_, state[118]);
    xor _4069_(_1740_, round_key[118], state[118]);
    and _4070_(_1741_, _1740_, _0779_);
    and _4071_(_1742_, _1741_, encrypting);
    and _4072_(_1743_, _1742_, _0781_);
    and _4073_(_1744_, _0799_, plaintext[118]);
    or _4074_(_1745_, _1744_, _1743_);
    and _4075_(_1746_, _1745_, _0794_);
    or _4076_(_0509_, _1746_, _1739_);
    and _4077_(_1747_, _0792_, state[119]);
    xor _4078_(_1748_, round_key[119], state[119]);
    and _4079_(_1749_, _1748_, _0779_);
    and _4080_(_1750_, _1749_, encrypting);
    and _4081_(_1751_, _1750_, _0781_);
    and _4082_(_1752_, _0799_, plaintext[119]);
    or _4083_(_1753_, _1752_, _1751_);
    and _4084_(_1754_, _1753_, _0794_);
    or _4085_(_0510_, _1754_, _1747_);
    and _4086_(_1755_, _0792_, state[120]);
    xor _4087_(_1756_, round_key[120], state[120]);
    and _4088_(_1757_, _1756_, _0779_);
    and _4089_(_1758_, _1757_, encrypting);
    and _4090_(_1759_, _1758_, _0781_);
    and _4091_(_1760_, _0799_, plaintext[120]);
    or _4092_(_1761_, _1760_, _1759_);
    and _4093_(_1762_, _1761_, _0794_);
    or _4094_(_0511_, _1762_, _1755_);
    and _4095_(_1763_, _0792_, state[121]);
    xor _4096_(_1764_, round_key[121], state[121]);
    and _4097_(_1765_, _1764_, _0779_);
    and _4098_(_1766_, _1765_, encrypting);
    and _4099_(_1767_, _1766_, _0781_);
    and _4100_(_1768_, _0799_, plaintext[121]);
    or _4101_(_1769_, _1768_, _1767_);
    and _4102_(_1770_, _1769_, _0794_);
    or _4103_(_0512_, _1770_, _1763_);
    and _4104_(_1771_, _0792_, state[122]);
    xor _4105_(_1772_, round_key[122], state[122]);
    and _4106_(_1773_, _1772_, _0779_);
    and _4107_(_1774_, _1773_, encrypting);
    and _4108_(_1775_, _1774_, _0781_);
    and _4109_(_1776_, _0799_, plaintext[122]);
    or _4110_(_1777_, _1776_, _1775_);
    and _4111_(_1778_, _1777_, _0794_);
    or _4112_(_0513_, _1778_, _1771_);
    and _4113_(_1779_, _0792_, state[123]);
    xor _4114_(_1780_, round_key[123], state[123]);
    and _4115_(_1781_, _1780_, _0779_);
    and _4116_(_1782_, _1781_, encrypting);
    and _4117_(_1783_, _1782_, _0781_);
    and _4118_(_1784_, _0799_, plaintext[123]);
    or _4119_(_1785_, _1784_, _1783_);
    and _4120_(_1786_, _1785_, _0794_);
    or _4121_(_0514_, _1786_, _1779_);
    and _4122_(_1787_, _0792_, state[124]);
    xor _4123_(_1788_, round_key[124], state[124]);
    and _4124_(_1789_, _1788_, _0779_);
    and _4125_(_1790_, _1789_, encrypting);
    and _4126_(_1791_, _1790_, _0781_);
    and _4127_(_1792_, _0799_, plaintext[124]);
    or _4128_(_1793_, _1792_, _1791_);
    and _4129_(_1794_, _1793_, _0794_);
    or _4130_(_0515_, _1794_, _1787_);
    and _4131_(_1795_, _0792_, state[125]);
    xor _4132_(_1796_, round_key[125], state[125]);
    and _4133_(_1797_, _1796_, _0779_);
    and _4134_(_1798_, _1797_, encrypting);
    and _4135_(_1799_, _1798_, _0781_);
    and _4136_(_1800_, _0799_, plaintext[125]);
    or _4137_(_1801_, _1800_, _1799_);
    and _4138_(_1802_, _1801_, _0794_);
    or _4139_(_0516_, _1802_, _1795_);
    and _4140_(_1803_, _0792_, state[126]);
    xor _4141_(_1804_, round_key[126], state[126]);
    and _4142_(_1805_, _1804_, _0779_);
    and _4143_(_1806_, _1805_, encrypting);
    and _4144_(_1807_, _1806_, _0781_);
    and _4145_(_1808_, _0799_, plaintext[126]);
    or _4146_(_1809_, _1808_, _1807_);
    and _4147_(_1810_, _1809_, _0794_);
    or _4148_(_0517_, _1810_, _1803_);
    and _4149_(_1811_, _0792_, state[127]);
    xor _4150_(_1812_, round_key[127], state[127]);
    and _4151_(_1813_, _1812_, _0779_);
    and _4152_(_1814_, _1813_, encrypting);
    and _4153_(_1815_, _1814_, _0781_);
    and _4154_(_1816_, _0799_, plaintext[127]);
    or _4155_(_1817_, _1816_, _1815_);
    and _4156_(_1818_, _1817_, _0794_);
    or _4157_(_0518_, _1818_, _1811_);
    and _4158_(_1819_, _0792_, round_key[0]);
    and _4159_(_1820_, _0779_, round_key[120]);
    and _4160_(_1821_, _1820_, encrypting);
    and _4161_(_1822_, _1821_, _0781_);
    and _4162_(_1823_, _0799_, cipher_key[0]);
    or _4163_(_1824_, _1823_, _1822_);
    and _4164_(_1825_, _1824_, _0794_);
    or _4165_(_0519_, _1825_, _1819_);
    and _4166_(_1826_, _0792_, round_key[1]);
    and _4167_(_1827_, _0779_, round_key[121]);
    and _4168_(_1828_, _1827_, encrypting);
    and _4169_(_1829_, _1828_, _0781_);
    and _4170_(_1830_, _0799_, cipher_key[1]);
    or _4171_(_1831_, _1830_, _1829_);
    and _4172_(_1832_, _1831_, _0794_);
    or _4173_(_0520_, _1832_, _1826_);
    and _4174_(_1833_, _0792_, round_key[2]);
    and _4175_(_1834_, _0779_, round_key[122]);
    and _4176_(_1835_, _1834_, encrypting);
    and _4177_(_1836_, _1835_, _0781_);
    and _4178_(_1837_, _0799_, cipher_key[2]);
    or _4179_(_1838_, _1837_, _1836_);
    and _4180_(_1839_, _1838_, _0794_);
    or _4181_(_0521_, _1839_, _1833_);
    and _4182_(_1840_, _0792_, round_key[3]);
    and _4183_(_1841_, _0779_, round_key[123]);
    and _4184_(_1842_, _1841_, encrypting);
    and _4185_(_1843_, _1842_, _0781_);
    and _4186_(_1844_, _0799_, cipher_key[3]);
    or _4187_(_1845_, _1844_, _1843_);
    and _4188_(_1846_, _1845_, _0794_);
    or _4189_(_0522_, _1846_, _1840_);
    and _4190_(_1847_, _0792_, round_key[4]);
    and _4191_(_1848_, _0779_, round_key[124]);
    and _4192_(_1849_, _1848_, encrypting);
    and _4193_(_1850_, _1849_, _0781_);
    and _4194_(_1851_, _0799_, cipher_key[4]);
    or _4195_(_1852_, _1851_, _1850_);
    and _4196_(_1853_, _1852_, _0794_);
    or _4197_(_0523_, _1853_, _1847_);
    and _4198_(_1854_, _0792_, round_key[5]);
    and _4199_(_1855_, _0779_, round_key[125]);
    and _4200_(_1856_, _1855_, encrypting);
    and _4201_(_1857_, _1856_, _0781_);
    and _4202_(_1858_, _0799_, cipher_key[5]);
    or _4203_(_1859_, _1858_, _1857_);
    and _4204_(_1860_, _1859_, _0794_);
    or _4205_(_0524_, _1860_, _1854_);
    and _4206_(_1861_, _0792_, round_key[6]);
    and _4207_(_1862_, _0779_, round_key[126]);
    and _4208_(_1863_, _1862_, encrypting);
    and _4209_(_1864_, _1863_, _0781_);
    and _4210_(_1865_, _0799_, cipher_key[6]);
    or _4211_(_1866_, _1865_, _1864_);
    and _4212_(_1867_, _1866_, _0794_);
    or _4213_(_0525_, _1867_, _1861_);
    and _4214_(_1868_, _0792_, round_key[7]);
    and _4215_(_1869_, _0779_, round_key[127]);
    and _4216_(_1870_, _1869_, encrypting);
    and _4217_(_1871_, _1870_, _0781_);
    and _4218_(_1872_, _0799_, cipher_key[7]);
    or _4219_(_1873_, _1872_, _1871_);
    and _4220_(_1874_, _1873_, _0794_);
    or _4221_(_0526_, _1874_, _1868_);
    and _4222_(_1875_, _0792_, round_key[8]);
    and _4223_(_1876_, _0779_, round_key[0]);
    and _4224_(_1877_, _1876_, encrypting);
    and _4225_(_1878_, _1877_, _0781_);
    and _4226_(_1879_, _0799_, cipher_key[8]);
    or _4227_(_1880_, _1879_, _1878_);
    and _4228_(_1881_, _1880_, _0794_);
    or _4229_(_0527_, _1881_, _1875_);
    and _4230_(_1882_, _0792_, round_key[9]);
    and _4231_(_1883_, _0779_, round_key[1]);
    and _4232_(_1884_, _1883_, encrypting);
    and _4233_(_1885_, _1884_, _0781_);
    and _4234_(_1886_, _0799_, cipher_key[9]);
    or _4235_(_1887_, _1886_, _1885_);
    and _4236_(_1888_, _1887_, _0794_);
    or _4237_(_0528_, _1888_, _1882_);
    and _4238_(_1889_, _0792_, round_key[10]);
    and _4239_(_1890_, _0779_, round_key[2]);
    and _4240_(_1891_, _1890_, encrypting);
    and _4241_(_1892_, _1891_, _0781_);
    and _4242_(_1893_, _0799_, cipher_key[10]);
    or _4243_(_1894_, _1893_, _1892_);
    and _4244_(_1895_, _1894_, _0794_);
    or _4245_(_0529_, _1895_, _1889_);
    and _4246_(_1896_, _0792_, round_key[11]);
    and _4247_(_1897_, _0779_, round_key[3]);
    and _4248_(_1898_, _1897_, encrypting);
    and _4249_(_1899_, _1898_, _0781_);
    and _4250_(_1900_, _0799_, cipher_key[11]);
    or _4251_(_1901_, _1900_, _1899_);
    and _4252_(_1902_, _1901_, _0794_);
    or _4253_(_0530_, _1902_, _1896_);
    and _4254_(_1903_, _0792_, round_key[12]);
    and _4255_(_1904_, _0779_, round_key[4]);
    and _4256_(_1905_, _1904_, encrypting);
    and _4257_(_1906_, _1905_, _0781_);
    and _4258_(_1907_, _0799_, cipher_key[12]);
    or _4259_(_1908_, _1907_, _1906_);
    and _4260_(_1909_, _1908_, _0794_);
    or _4261_(_0531_, _1909_, _1903_);
    and _4262_(_1910_, _0792_, round_key[13]);
    and _4263_(_1911_, _0779_, round_key[5]);
    and _4264_(_1912_, _1911_, encrypting);
    and _4265_(_1913_, _1912_, _0781_);
    and _4266_(_1914_, _0799_, cipher_key[13]);
    or _4267_(_1915_, _1914_, _1913_);
    and _4268_(_1916_, _1915_, _0794_);
    or _4269_(_0532_, _1916_, _1910_);
    and _4270_(_1917_, _0792_, round_key[14]);
    and _4271_(_1918_, _0779_, round_key[6]);
    and _4272_(_1919_, _1918_, encrypting);
    and _4273_(_1920_, _1919_, _0781_);
    and _4274_(_1921_, _0799_, cipher_key[14]);
    or _4275_(_1922_, _1921_, _1920_);
    and _4276_(_1923_, _1922_, _0794_);
    or _4277_(_0533_, _1923_, _1917_);
    and _4278_(_1924_, _0792_, round_key[15]);
    and _4279_(_1925_, _0779_, round_key[7]);
    and _4280_(_1926_, _1925_, encrypting);
    and _4281_(_1927_, _1926_, _0781_);
    and _4282_(_1928_, _0799_, cipher_key[15]);
    or _4283_(_1929_, _1928_, _1927_);
    and _4284_(_1930_, _1929_, _0794_);
    or _4285_(_0534_, _1930_, _1924_);
    and _4286_(_1931_, _0792_, round_key[16]);
    and _4287_(_1932_, _0779_, round_key[8]);
    and _4288_(_1933_, _1932_, encrypting);
    and _4289_(_1934_, _1933_, _0781_);
    and _4290_(_1935_, _0799_, cipher_key[16]);
    or _4291_(_1936_, _1935_, _1934_);
    and _4292_(_1937_, _1936_, _0794_);
    or _4293_(_0535_, _1937_, _1931_);
    and _4294_(_1938_, _0792_, round_key[17]);
    and _4295_(_1939_, _0779_, round_key[9]);
    and _4296_(_1940_, _1939_, encrypting);
    and _4297_(_1941_, _1940_, _0781_);
    and _4298_(_1942_, _0799_, cipher_key[17]);
    or _4299_(_1943_, _1942_, _1941_);
    and _4300_(_1944_, _1943_, _0794_);
    or _4301_(_0536_, _1944_, _1938_);
    and _4302_(_1945_, _0792_, round_key[18]);
    and _4303_(_1946_, _0779_, round_key[10]);
    and _4304_(_1947_, _1946_, encrypting);
    and _4305_(_1948_, _1947_, _0781_);
    and _4306_(_1949_, _0799_, cipher_key[18]);
    or _4307_(_1950_, _1949_, _1948_);
    and _4308_(_1951_, _1950_, _0794_);
    or _4309_(_0537_, _1951_, _1945_);
    and _4310_(_1952_, _0792_, round_key[19]);
    and _4311_(_1953_, _0779_, round_key[11]);
    and _4312_(_1954_, _1953_, encrypting);
    and _4313_(_1955_, _1954_, _0781_);
    and _4314_(_1956_, _0799_, cipher_key[19]);
    or _4315_(_1957_, _1956_, _1955_);
    and _4316_(_1958_, _1957_, _0794_);
    or _4317_(_0538_, _1958_, _1952_);
    and _4318_(_1959_, _0792_, round_key[20]);
    and _4319_(_1960_, _0779_, round_key[12]);
    and _4320_(_1961_, _1960_, encrypting);
    and _4321_(_1962_, _1961_, _0781_);
    and _4322_(_1963_, _0799_, cipher_key[20]);
    or _4323_(_1964_, _1963_, _1962_);
    and _4324_(_1965_, _1964_, _0794_);
    or _4325_(_0539_, _1965_, _1959_);
    and _4326_(_1966_, _0792_, round_key[21]);
    and _4327_(_1967_, _0779_, round_key[13]);
    and _4328_(_1968_, _1967_, encrypting);
    and _4329_(_1969_, _1968_, _0781_);
    and _4330_(_1970_, _0799_, cipher_key[21]);
    or _4331_(_1971_, _1970_, _1969_);
    and _4332_(_1972_, _1971_, _0794_);
    or _4333_(_0540_, _1972_, _1966_);
    and _4334_(_1973_, _0792_, round_key[22]);
    and _4335_(_1974_, _0779_, round_key[14]);
    and _4336_(_1975_, _1974_, encrypting);
    and _4337_(_1976_, _1975_, _0781_);
    and _4338_(_1977_, _0799_, cipher_key[22]);
    or _4339_(_1978_, _1977_, _1976_);
    and _4340_(_1979_, _1978_, _0794_);
    or _4341_(_0541_, _1979_, _1973_);
    and _4342_(_1980_, _0792_, round_key[23]);
    and _4343_(_1981_, _0779_, round_key[15]);
    and _4344_(_1982_, _1981_, encrypting);
    and _4345_(_1983_, _1982_, _0781_);
    and _4346_(_1984_, _0799_, cipher_key[23]);
    or _4347_(_1985_, _1984_, _1983_);
    and _4348_(_1986_, _1985_, _0794_);
    or _4349_(_0542_, _1986_, _1980_);
    and _4350_(_1987_, _0792_, round_key[24]);
    and _4351_(_1988_, _0779_, round_key[16]);
    and _4352_(_1989_, _1988_, encrypting);
    and _4353_(_1990_, _1989_, _0781_);
    and _4354_(_1991_, _0799_, cipher_key[24]);
    or _4355_(_1992_, _1991_, _1990_);
    and _4356_(_1993_, _1992_, _0794_);
    or _4357_(_0543_, _1993_, _1987_);
    and _4358_(_1994_, _0792_, round_key[25]);
    and _4359_(_1995_, _0779_, round_key[17]);
    and _4360_(_1996_, _1995_, encrypting);
    and _4361_(_1997_, _1996_, _0781_);
    and _4362_(_1998_, _0799_, cipher_key[25]);
    or _4363_(_1999_, _1998_, _1997_);
    and _4364_(_2000_, _1999_, _0794_);
    or _4365_(_0544_, _2000_, _1994_);
    and _4366_(_2001_, _0792_, round_key[26]);
    and _4367_(_2002_, _0779_, round_key[18]);
    and _4368_(_2003_, _2002_, encrypting);
    and _4369_(_2004_, _2003_, _0781_);
    and _4370_(_2005_, _0799_, cipher_key[26]);
    or _4371_(_2006_, _2005_, _2004_);
    and _4372_(_2007_, _2006_, _0794_);
    or _4373_(_0545_, _2007_, _2001_);
    and _4374_(_2008_, _0792_, round_key[27]);
    and _4375_(_2009_, _0779_, round_key[19]);
    and _4376_(_2010_, _2009_, encrypting);
    and _4377_(_2011_, _2010_, _0781_);
    and _4378_(_2012_, _0799_, cipher_key[27]);
    or _4379_(_2013_, _2012_, _2011_);
    and _4380_(_2014_, _2013_, _0794_);
    or _4381_(_0546_, _2014_, _2008_);
    and _4382_(_2015_, _0792_, round_key[28]);
    and _4383_(_2016_, _0779_, round_key[20]);
    and _4384_(_2017_, _2016_, encrypting);
    and _4385_(_2018_, _2017_, _0781_);
    and _4386_(_2019_, _0799_, cipher_key[28]);
    or _4387_(_2020_, _2019_, _2018_);
    and _4388_(_2021_, _2020_, _0794_);
    or _4389_(_0547_, _2021_, _2015_);
    and _4390_(_2022_, _0792_, round_key[29]);
    and _4391_(_2023_, _0779_, round_key[21]);
    and _4392_(_2024_, _2023_, encrypting);
    and _4393_(_2025_, _2024_, _0781_);
    and _4394_(_2026_, _0799_, cipher_key[29]);
    or _4395_(_2027_, _2026_, _2025_);
    and _4396_(_2028_, _2027_, _0794_);
    or _4397_(_0548_, _2028_, _2022_);
    and _4398_(_2029_, _0792_, round_key[30]);
    and _4399_(_2030_, _0779_, round_key[22]);
    and _4400_(_2031_, _2030_, encrypting);
    and _4401_(_2032_, _2031_, _0781_);
    and _4402_(_2033_, _0799_, cipher_key[30]);
    or _4403_(_2034_, _2033_, _2032_);
    and _4404_(_2035_, _2034_, _0794_);
    or _4405_(_0549_, _2035_, _2029_);
    and _4406_(_2036_, _0792_, round_key[31]);
    and _4407_(_2037_, _0779_, round_key[23]);
    and _4408_(_2038_, _2037_, encrypting);
    and _4409_(_2039_, _2038_, _0781_);
    and _4410_(_2040_, _0799_, cipher_key[31]);
    or _4411_(_2041_, _2040_, _2039_);
    and _4412_(_2042_, _2041_, _0794_);
    or _4413_(_0550_, _2042_, _2036_);
    and _4414_(_2043_, _0792_, round_key[32]);
    and _4415_(_2044_, _0779_, round_key[24]);
    and _4416_(_2045_, _2044_, encrypting);
    and _4417_(_2046_, _2045_, _0781_);
    and _4418_(_2047_, _0799_, cipher_key[32]);
    or _4419_(_2048_, _2047_, _2046_);
    and _4420_(_2049_, _2048_, _0794_);
    or _4421_(_0551_, _2049_, _2043_);
    and _4422_(_2050_, _0792_, round_key[33]);
    and _4423_(_2051_, _0779_, round_key[25]);
    and _4424_(_2052_, _2051_, encrypting);
    and _4425_(_2053_, _2052_, _0781_);
    and _4426_(_2054_, _0799_, cipher_key[33]);
    or _4427_(_2055_, _2054_, _2053_);
    and _4428_(_2056_, _2055_, _0794_);
    or _4429_(_0552_, _2056_, _2050_);
    and _4430_(_2057_, _0792_, round_key[34]);
    and _4431_(_2058_, _0779_, round_key[26]);
    and _4432_(_2059_, _2058_, encrypting);
    and _4433_(_2060_, _2059_, _0781_);
    and _4434_(_2061_, _0799_, cipher_key[34]);
    or _4435_(_2062_, _2061_, _2060_);
    and _4436_(_2063_, _2062_, _0794_);
    or _4437_(_0553_, _2063_, _2057_);
    and _4438_(_2064_, _0792_, round_key[35]);
    and _4439_(_2065_, _0779_, round_key[27]);
    and _4440_(_2066_, _2065_, encrypting);
    and _4441_(_2067_, _2066_, _0781_);
    and _4442_(_2068_, _0799_, cipher_key[35]);
    or _4443_(_2069_, _2068_, _2067_);
    and _4444_(_2070_, _2069_, _0794_);
    or _4445_(_0554_, _2070_, _2064_);
    and _4446_(_2071_, _0792_, round_key[36]);
    and _4447_(_2072_, _0779_, round_key[28]);
    and _4448_(_2073_, _2072_, encrypting);
    and _4449_(_2074_, _2073_, _0781_);
    and _4450_(_2075_, _0799_, cipher_key[36]);
    or _4451_(_2076_, _2075_, _2074_);
    and _4452_(_2077_, _2076_, _0794_);
    or _4453_(_0555_, _2077_, _2071_);
    and _4454_(_2078_, _0792_, round_key[37]);
    and _4455_(_2079_, _0779_, round_key[29]);
    and _4456_(_2080_, _2079_, encrypting);
    and _4457_(_2081_, _2080_, _0781_);
    and _4458_(_2082_, _0799_, cipher_key[37]);
    or _4459_(_2083_, _2082_, _2081_);
    and _4460_(_2084_, _2083_, _0794_);
    or _4461_(_0556_, _2084_, _2078_);
    and _4462_(_2085_, _0792_, round_key[38]);
    and _4463_(_2086_, _0779_, round_key[30]);
    and _4464_(_2087_, _2086_, encrypting);
    and _4465_(_2088_, _2087_, _0781_);
    and _4466_(_2089_, _0799_, cipher_key[38]);
    or _4467_(_2090_, _2089_, _2088_);
    and _4468_(_2091_, _2090_, _0794_);
    or _4469_(_0557_, _2091_, _2085_);
    and _4470_(_2092_, _0792_, round_key[39]);
    and _4471_(_2093_, _0779_, round_key[31]);
    and _4472_(_2094_, _2093_, encrypting);
    and _4473_(_2095_, _2094_, _0781_);
    and _4474_(_2096_, _0799_, cipher_key[39]);
    or _4475_(_2097_, _2096_, _2095_);
    and _4476_(_2098_, _2097_, _0794_);
    or _4477_(_0558_, _2098_, _2092_);
    and _4478_(_2099_, _0792_, round_key[40]);
    and _4479_(_2100_, _0779_, round_key[32]);
    and _4480_(_2101_, _2100_, encrypting);
    and _4481_(_2102_, _2101_, _0781_);
    and _4482_(_2103_, _0799_, cipher_key[40]);
    or _4483_(_2104_, _2103_, _2102_);
    and _4484_(_2105_, _2104_, _0794_);
    or _4485_(_0559_, _2105_, _2099_);
    and _4486_(_2106_, _0792_, round_key[41]);
    and _4487_(_2107_, _0779_, round_key[33]);
    and _4488_(_2108_, _2107_, encrypting);
    and _4489_(_2109_, _2108_, _0781_);
    and _4490_(_2110_, _0799_, cipher_key[41]);
    or _4491_(_2111_, _2110_, _2109_);
    and _4492_(_2112_, _2111_, _0794_);
    or _4493_(_0560_, _2112_, _2106_);
    and _4494_(_2113_, _0792_, round_key[42]);
    and _4495_(_2114_, _0779_, round_key[34]);
    and _4496_(_2115_, _2114_, encrypting);
    and _4497_(_2116_, _2115_, _0781_);
    and _4498_(_2117_, _0799_, cipher_key[42]);
    or _4499_(_2118_, _2117_, _2116_);
    and _4500_(_2119_, _2118_, _0794_);
    or _4501_(_0561_, _2119_, _2113_);
    and _4502_(_2120_, _0792_, round_key[43]);
    and _4503_(_2121_, _0779_, round_key[35]);
    and _4504_(_2122_, _2121_, encrypting);
    and _4505_(_2123_, _2122_, _0781_);
    and _4506_(_2124_, _0799_, cipher_key[43]);
    or _4507_(_2125_, _2124_, _2123_);
    and _4508_(_2126_, _2125_, _0794_);
    or _4509_(_0562_, _2126_, _2120_);
    and _4510_(_2127_, _0792_, round_key[44]);
    and _4511_(_2128_, _0779_, round_key[36]);
    and _4512_(_2129_, _2128_, encrypting);
    and _4513_(_2130_, _2129_, _0781_);
    and _4514_(_2131_, _0799_, cipher_key[44]);
    or _4515_(_2132_, _2131_, _2130_);
    and _4516_(_2133_, _2132_, _0794_);
    or _4517_(_0563_, _2133_, _2127_);
    and _4518_(_2134_, _0792_, round_key[45]);
    and _4519_(_2135_, _0779_, round_key[37]);
    and _4520_(_2136_, _2135_, encrypting);
    and _4521_(_2137_, _2136_, _0781_);
    and _4522_(_2138_, _0799_, cipher_key[45]);
    or _4523_(_2139_, _2138_, _2137_);
    and _4524_(_2140_, _2139_, _0794_);
    or _4525_(_0564_, _2140_, _2134_);
    and _4526_(_2141_, _0792_, round_key[46]);
    and _4527_(_2142_, _0779_, round_key[38]);
    and _4528_(_2143_, _2142_, encrypting);
    and _4529_(_2144_, _2143_, _0781_);
    and _4530_(_2145_, _0799_, cipher_key[46]);
    or _4531_(_2146_, _2145_, _2144_);
    and _4532_(_2147_, _2146_, _0794_);
    or _4533_(_0565_, _2147_, _2141_);
    and _4534_(_2148_, _0792_, round_key[47]);
    and _4535_(_2149_, _0779_, round_key[39]);
    and _4536_(_2150_, _2149_, encrypting);
    and _4537_(_2151_, _2150_, _0781_);
    and _4538_(_2152_, _0799_, cipher_key[47]);
    or _4539_(_2153_, _2152_, _2151_);
    and _4540_(_2154_, _2153_, _0794_);
    or _4541_(_0566_, _2154_, _2148_);
    and _4542_(_2155_, _0792_, round_key[48]);
    and _4543_(_2156_, _0779_, round_key[40]);
    and _4544_(_2157_, _2156_, encrypting);
    and _4545_(_2158_, _2157_, _0781_);
    and _4546_(_2159_, _0799_, cipher_key[48]);
    or _4547_(_2160_, _2159_, _2158_);
    and _4548_(_2161_, _2160_, _0794_);
    or _4549_(_0567_, _2161_, _2155_);
    and _4550_(_2162_, _0792_, round_key[49]);
    and _4551_(_2163_, _0779_, round_key[41]);
    and _4552_(_2164_, _2163_, encrypting);
    and _4553_(_2165_, _2164_, _0781_);
    and _4554_(_2166_, _0799_, cipher_key[49]);
    or _4555_(_2167_, _2166_, _2165_);
    and _4556_(_2168_, _2167_, _0794_);
    or _4557_(_0568_, _2168_, _2162_);
    and _4558_(_2169_, _0792_, round_key[50]);
    and _4559_(_2170_, _0779_, round_key[42]);
    and _4560_(_2171_, _2170_, encrypting);
    and _4561_(_2172_, _2171_, _0781_);
    and _4562_(_2173_, _0799_, cipher_key[50]);
    or _4563_(_2174_, _2173_, _2172_);
    and _4564_(_2175_, _2174_, _0794_);
    or _4565_(_0569_, _2175_, _2169_);
    and _4566_(_2176_, _0792_, round_key[51]);
    and _4567_(_2177_, _0779_, round_key[43]);
    and _4568_(_2178_, _2177_, encrypting);
    and _4569_(_2179_, _2178_, _0781_);
    and _4570_(_2180_, _0799_, cipher_key[51]);
    or _4571_(_2181_, _2180_, _2179_);
    and _4572_(_2182_, _2181_, _0794_);
    or _4573_(_0570_, _2182_, _2176_);
    and _4574_(_2183_, _0792_, round_key[52]);
    and _4575_(_2184_, _0779_, round_key[44]);
    and _4576_(_2185_, _2184_, encrypting);
    and _4577_(_2186_, _2185_, _0781_);
    and _4578_(_2187_, _0799_, cipher_key[52]);
    or _4579_(_2188_, _2187_, _2186_);
    and _4580_(_2189_, _2188_, _0794_);
    or _4581_(_0571_, _2189_, _2183_);
    and _4582_(_2190_, _0792_, round_key[53]);
    and _4583_(_2191_, _0779_, round_key[45]);
    and _4584_(_2192_, _2191_, encrypting);
    and _4585_(_2193_, _2192_, _0781_);
    and _4586_(_2194_, _0799_, cipher_key[53]);
    or _4587_(_2195_, _2194_, _2193_);
    and _4588_(_2196_, _2195_, _0794_);
    or _4589_(_0572_, _2196_, _2190_);
    and _4590_(_2197_, _0792_, round_key[54]);
    and _4591_(_2198_, _0779_, round_key[46]);
    and _4592_(_2199_, _2198_, encrypting);
    and _4593_(_2200_, _2199_, _0781_);
    and _4594_(_2201_, _0799_, cipher_key[54]);
    or _4595_(_2202_, _2201_, _2200_);
    and _4596_(_2203_, _2202_, _0794_);
    or _4597_(_0573_, _2203_, _2197_);
    and _4598_(_2204_, _0792_, round_key[55]);
    and _4599_(_2205_, _0779_, round_key[47]);
    and _4600_(_2206_, _2205_, encrypting);
    and _4601_(_2207_, _2206_, _0781_);
    and _4602_(_2208_, _0799_, cipher_key[55]);
    or _4603_(_2209_, _2208_, _2207_);
    and _4604_(_2210_, _2209_, _0794_);
    or _4605_(_0574_, _2210_, _2204_);
    and _4606_(_2211_, _0792_, round_key[56]);
    and _4607_(_2212_, _0779_, round_key[48]);
    and _4608_(_2213_, _2212_, encrypting);
    and _4609_(_2214_, _2213_, _0781_);
    and _4610_(_2215_, _0799_, cipher_key[56]);
    or _4611_(_2216_, _2215_, _2214_);
    and _4612_(_2217_, _2216_, _0794_);
    or _4613_(_0575_, _2217_, _2211_);
    and _4614_(_2218_, _0792_, round_key[57]);
    and _4615_(_2219_, _0779_, round_key[49]);
    and _4616_(_2220_, _2219_, encrypting);
    and _4617_(_2221_, _2220_, _0781_);
    and _4618_(_2222_, _0799_, cipher_key[57]);
    or _4619_(_2223_, _2222_, _2221_);
    and _4620_(_2224_, _2223_, _0794_);
    or _4621_(_0576_, _2224_, _2218_);
    and _4622_(_2225_, _0792_, round_key[58]);
    and _4623_(_2226_, _0779_, round_key[50]);
    and _4624_(_2227_, _2226_, encrypting);
    and _4625_(_2228_, _2227_, _0781_);
    and _4626_(_2229_, _0799_, cipher_key[58]);
    or _4627_(_2230_, _2229_, _2228_);
    and _4628_(_2231_, _2230_, _0794_);
    or _4629_(_0577_, _2231_, _2225_);
    and _4630_(_2232_, _0792_, round_key[59]);
    and _4631_(_2233_, _0779_, round_key[51]);
    and _4632_(_2234_, _2233_, encrypting);
    and _4633_(_2235_, _2234_, _0781_);
    and _4634_(_2236_, _0799_, cipher_key[59]);
    or _4635_(_2237_, _2236_, _2235_);
    and _4636_(_2238_, _2237_, _0794_);
    or _4637_(_0578_, _2238_, _2232_);
    and _4638_(_2239_, _0792_, round_key[60]);
    and _4639_(_2240_, _0779_, round_key[52]);
    and _4640_(_2241_, _2240_, encrypting);
    and _4641_(_2242_, _2241_, _0781_);
    and _4642_(_2243_, _0799_, cipher_key[60]);
    or _4643_(_2244_, _2243_, _2242_);
    and _4644_(_2245_, _2244_, _0794_);
    or _4645_(_0579_, _2245_, _2239_);
    and _4646_(_2246_, _0792_, round_key[61]);
    and _4647_(_2247_, _0779_, round_key[53]);
    and _4648_(_2248_, _2247_, encrypting);
    and _4649_(_2249_, _2248_, _0781_);
    and _4650_(_2250_, _0799_, cipher_key[61]);
    or _4651_(_2251_, _2250_, _2249_);
    and _4652_(_2252_, _2251_, _0794_);
    or _4653_(_0580_, _2252_, _2246_);
    and _4654_(_2253_, _0792_, round_key[62]);
    and _4655_(_2254_, _0779_, round_key[54]);
    and _4656_(_2255_, _2254_, encrypting);
    and _4657_(_2256_, _2255_, _0781_);
    and _4658_(_2257_, _0799_, cipher_key[62]);
    or _4659_(_2258_, _2257_, _2256_);
    and _4660_(_2259_, _2258_, _0794_);
    or _4661_(_0581_, _2259_, _2253_);
    and _4662_(_2260_, _0792_, round_key[63]);
    and _4663_(_2261_, _0779_, round_key[55]);
    and _4664_(_2262_, _2261_, encrypting);
    and _4665_(_2263_, _2262_, _0781_);
    and _4666_(_2264_, _0799_, cipher_key[63]);
    or _4667_(_2265_, _2264_, _2263_);
    and _4668_(_2266_, _2265_, _0794_);
    or _4669_(_0582_, _2266_, _2260_);
    and _4670_(_2267_, _0792_, round_key[64]);
    and _4671_(_2268_, _0779_, round_key[56]);
    and _4672_(_2269_, _2268_, encrypting);
    and _4673_(_2270_, _2269_, _0781_);
    and _4674_(_2271_, _0799_, cipher_key[64]);
    or _4675_(_2272_, _2271_, _2270_);
    and _4676_(_2273_, _2272_, _0794_);
    or _4677_(_0583_, _2273_, _2267_);
    and _4678_(_2274_, _0792_, round_key[65]);
    and _4679_(_2275_, _0779_, round_key[57]);
    and _4680_(_2276_, _2275_, encrypting);
    and _4681_(_2277_, _2276_, _0781_);
    and _4682_(_2278_, _0799_, cipher_key[65]);
    or _4683_(_2279_, _2278_, _2277_);
    and _4684_(_2280_, _2279_, _0794_);
    or _4685_(_0584_, _2280_, _2274_);
    and _4686_(_2281_, _0792_, round_key[66]);
    and _4687_(_2282_, _0779_, round_key[58]);
    and _4688_(_2283_, _2282_, encrypting);
    and _4689_(_2284_, _2283_, _0781_);
    and _4690_(_2285_, _0799_, cipher_key[66]);
    or _4691_(_2286_, _2285_, _2284_);
    and _4692_(_2287_, _2286_, _0794_);
    or _4693_(_0585_, _2287_, _2281_);
    and _4694_(_2288_, _0792_, round_key[67]);
    and _4695_(_2289_, _0779_, round_key[59]);
    and _4696_(_2290_, _2289_, encrypting);
    and _4697_(_2291_, _2290_, _0781_);
    and _4698_(_2292_, _0799_, cipher_key[67]);
    or _4699_(_2293_, _2292_, _2291_);
    and _4700_(_2294_, _2293_, _0794_);
    or _4701_(_0586_, _2294_, _2288_);
    and _4702_(_2295_, _0792_, round_key[68]);
    and _4703_(_2296_, _0779_, round_key[60]);
    and _4704_(_2297_, _2296_, encrypting);
    and _4705_(_2298_, _2297_, _0781_);
    and _4706_(_2299_, _0799_, cipher_key[68]);
    or _4707_(_2300_, _2299_, _2298_);
    and _4708_(_2301_, _2300_, _0794_);
    or _4709_(_0587_, _2301_, _2295_);
    and _4710_(_2302_, _0792_, round_key[69]);
    and _4711_(_2303_, _0779_, round_key[61]);
    and _4712_(_2304_, _2303_, encrypting);
    and _4713_(_2305_, _2304_, _0781_);
    and _4714_(_2306_, _0799_, cipher_key[69]);
    or _4715_(_2307_, _2306_, _2305_);
    and _4716_(_2308_, _2307_, _0794_);
    or _4717_(_0588_, _2308_, _2302_);
    and _4718_(_2309_, _0792_, round_key[70]);
    and _4719_(_2310_, _0779_, round_key[62]);
    and _4720_(_2311_, _2310_, encrypting);
    and _4721_(_2312_, _2311_, _0781_);
    and _4722_(_2313_, _0799_, cipher_key[70]);
    or _4723_(_2314_, _2313_, _2312_);
    and _4724_(_2315_, _2314_, _0794_);
    or _4725_(_0589_, _2315_, _2309_);
    and _4726_(_2316_, _0792_, round_key[71]);
    and _4727_(_2317_, _0779_, round_key[63]);
    and _4728_(_2318_, _2317_, encrypting);
    and _4729_(_2319_, _2318_, _0781_);
    and _4730_(_2320_, _0799_, cipher_key[71]);
    or _4731_(_2321_, _2320_, _2319_);
    and _4732_(_2322_, _2321_, _0794_);
    or _4733_(_0590_, _2322_, _2316_);
    and _4734_(_2323_, _0792_, round_key[72]);
    and _4735_(_2324_, _0779_, round_key[64]);
    and _4736_(_2325_, _2324_, encrypting);
    and _4737_(_2326_, _2325_, _0781_);
    and _4738_(_2327_, _0799_, cipher_key[72]);
    or _4739_(_2328_, _2327_, _2326_);
    and _4740_(_2329_, _2328_, _0794_);
    or _4741_(_0591_, _2329_, _2323_);
    and _4742_(_2330_, _0792_, round_key[73]);
    and _4743_(_2331_, _0779_, round_key[65]);
    and _4744_(_2332_, _2331_, encrypting);
    and _4745_(_2333_, _2332_, _0781_);
    and _4746_(_2334_, _0799_, cipher_key[73]);
    or _4747_(_2335_, _2334_, _2333_);
    and _4748_(_2336_, _2335_, _0794_);
    or _4749_(_0592_, _2336_, _2330_);
    and _4750_(_2337_, _0792_, round_key[74]);
    and _4751_(_2338_, _0779_, round_key[66]);
    and _4752_(_2339_, _2338_, encrypting);
    and _4753_(_2340_, _2339_, _0781_);
    and _4754_(_2341_, _0799_, cipher_key[74]);
    or _4755_(_2342_, _2341_, _2340_);
    and _4756_(_2343_, _2342_, _0794_);
    or _4757_(_0593_, _2343_, _2337_);
    and _4758_(_2344_, _0792_, round_key[75]);
    and _4759_(_2345_, _0779_, round_key[67]);
    and _4760_(_2346_, _2345_, encrypting);
    and _4761_(_2347_, _2346_, _0781_);
    and _4762_(_2348_, _0799_, cipher_key[75]);
    or _4763_(_2349_, _2348_, _2347_);
    and _4764_(_2350_, _2349_, _0794_);
    or _4765_(_0594_, _2350_, _2344_);
    and _4766_(_2351_, _0792_, round_key[76]);
    and _4767_(_2352_, _0779_, round_key[68]);
    and _4768_(_2353_, _2352_, encrypting);
    and _4769_(_2354_, _2353_, _0781_);
    and _4770_(_2355_, _0799_, cipher_key[76]);
    or _4771_(_2356_, _2355_, _2354_);
    and _4772_(_2357_, _2356_, _0794_);
    or _4773_(_0595_, _2357_, _2351_);
    and _4774_(_2358_, _0792_, round_key[77]);
    and _4775_(_2359_, _0779_, round_key[69]);
    and _4776_(_2360_, _2359_, encrypting);
    and _4777_(_2361_, _2360_, _0781_);
    and _4778_(_2362_, _0799_, cipher_key[77]);
    or _4779_(_2363_, _2362_, _2361_);
    and _4780_(_2364_, _2363_, _0794_);
    or _4781_(_0596_, _2364_, _2358_);
    and _4782_(_2365_, _0792_, round_key[78]);
    and _4783_(_2366_, _0779_, round_key[70]);
    and _4784_(_2367_, _2366_, encrypting);
    and _4785_(_2368_, _2367_, _0781_);
    and _4786_(_2369_, _0799_, cipher_key[78]);
    or _4787_(_2370_, _2369_, _2368_);
    and _4788_(_2371_, _2370_, _0794_);
    or _4789_(_0597_, _2371_, _2365_);
    and _4790_(_2372_, _0792_, round_key[79]);
    and _4791_(_2373_, _0779_, round_key[71]);
    and _4792_(_2374_, _2373_, encrypting);
    and _4793_(_2375_, _2374_, _0781_);
    and _4794_(_2376_, _0799_, cipher_key[79]);
    or _4795_(_2377_, _2376_, _2375_);
    and _4796_(_2378_, _2377_, _0794_);
    or _4797_(_0598_, _2378_, _2372_);
    and _4798_(_2379_, _0792_, round_key[80]);
    and _4799_(_2380_, _0779_, round_key[72]);
    and _4800_(_2381_, _2380_, encrypting);
    and _4801_(_2382_, _2381_, _0781_);
    and _4802_(_2383_, _0799_, cipher_key[80]);
    or _4803_(_2384_, _2383_, _2382_);
    and _4804_(_2385_, _2384_, _0794_);
    or _4805_(_0599_, _2385_, _2379_);
    and _4806_(_2386_, _0792_, round_key[81]);
    and _4807_(_2387_, _0779_, round_key[73]);
    and _4808_(_2388_, _2387_, encrypting);
    and _4809_(_2389_, _2388_, _0781_);
    and _4810_(_2390_, _0799_, cipher_key[81]);
    or _4811_(_2391_, _2390_, _2389_);
    and _4812_(_2392_, _2391_, _0794_);
    or _4813_(_0600_, _2392_, _2386_);
    and _4814_(_2393_, _0792_, round_key[82]);
    and _4815_(_2394_, _0779_, round_key[74]);
    and _4816_(_2395_, _2394_, encrypting);
    and _4817_(_2396_, _2395_, _0781_);
    and _4818_(_2397_, _0799_, cipher_key[82]);
    or _4819_(_2398_, _2397_, _2396_);
    and _4820_(_2399_, _2398_, _0794_);
    or _4821_(_0601_, _2399_, _2393_);
    and _4822_(_2400_, _0792_, round_key[83]);
    and _4823_(_2401_, _0779_, round_key[75]);
    and _4824_(_2402_, _2401_, encrypting);
    and _4825_(_2403_, _2402_, _0781_);
    and _4826_(_2404_, _0799_, cipher_key[83]);
    or _4827_(_2405_, _2404_, _2403_);
    and _4828_(_2406_, _2405_, _0794_);
    or _4829_(_0602_, _2406_, _2400_);
    and _4830_(_2407_, _0792_, round_key[84]);
    and _4831_(_2408_, _0779_, round_key[76]);
    and _4832_(_2409_, _2408_, encrypting);
    and _4833_(_2410_, _2409_, _0781_);
    and _4834_(_2411_, _0799_, cipher_key[84]);
    or _4835_(_2412_, _2411_, _2410_);
    and _4836_(_2413_, _2412_, _0794_);
    or _4837_(_0603_, _2413_, _2407_);
    and _4838_(_2414_, _0792_, round_key[85]);
    and _4839_(_2415_, _0779_, round_key[77]);
    and _4840_(_2416_, _2415_, encrypting);
    and _4841_(_2417_, _2416_, _0781_);
    and _4842_(_2418_, _0799_, cipher_key[85]);
    or _4843_(_2419_, _2418_, _2417_);
    and _4844_(_2420_, _2419_, _0794_);
    or _4845_(_0604_, _2420_, _2414_);
    and _4846_(_2421_, _0792_, round_key[86]);
    and _4847_(_2422_, _0779_, round_key[78]);
    and _4848_(_2423_, _2422_, encrypting);
    and _4849_(_2424_, _2423_, _0781_);
    and _4850_(_2425_, _0799_, cipher_key[86]);
    or _4851_(_2426_, _2425_, _2424_);
    and _4852_(_2427_, _2426_, _0794_);
    or _4853_(_0605_, _2427_, _2421_);
    and _4854_(_2428_, _0792_, round_key[87]);
    and _4855_(_2429_, _0779_, round_key[79]);
    and _4856_(_2430_, _2429_, encrypting);
    and _4857_(_2431_, _2430_, _0781_);
    and _4858_(_2432_, _0799_, cipher_key[87]);
    or _4859_(_2433_, _2432_, _2431_);
    and _4860_(_2434_, _2433_, _0794_);
    or _4861_(_0606_, _2434_, _2428_);
    and _4862_(_2435_, _0792_, round_key[88]);
    and _4863_(_2436_, _0779_, round_key[80]);
    and _4864_(_2437_, _2436_, encrypting);
    and _4865_(_2438_, _2437_, _0781_);
    and _4866_(_2439_, _0799_, cipher_key[88]);
    or _4867_(_2440_, _2439_, _2438_);
    and _4868_(_2441_, _2440_, _0794_);
    or _4869_(_0607_, _2441_, _2435_);
    and _4870_(_2442_, _0792_, round_key[89]);
    and _4871_(_2443_, _0779_, round_key[81]);
    and _4872_(_2444_, _2443_, encrypting);
    and _4873_(_2445_, _2444_, _0781_);
    and _4874_(_2446_, _0799_, cipher_key[89]);
    or _4875_(_2447_, _2446_, _2445_);
    and _4876_(_2448_, _2447_, _0794_);
    or _4877_(_0608_, _2448_, _2442_);
    and _4878_(_2449_, _0792_, round_key[90]);
    and _4879_(_2450_, _0779_, round_key[82]);
    and _4880_(_2451_, _2450_, encrypting);
    and _4881_(_2452_, _2451_, _0781_);
    and _4882_(_2453_, _0799_, cipher_key[90]);
    or _4883_(_2454_, _2453_, _2452_);
    and _4884_(_2455_, _2454_, _0794_);
    or _4885_(_0609_, _2455_, _2449_);
    and _4886_(_2456_, _0792_, round_key[91]);
    and _4887_(_2457_, _0779_, round_key[83]);
    and _4888_(_2458_, _2457_, encrypting);
    and _4889_(_2459_, _2458_, _0781_);
    and _4890_(_2460_, _0799_, cipher_key[91]);
    or _4891_(_2461_, _2460_, _2459_);
    and _4892_(_2462_, _2461_, _0794_);
    or _4893_(_0610_, _2462_, _2456_);
    and _4894_(_2463_, _0792_, round_key[92]);
    and _4895_(_2464_, _0779_, round_key[84]);
    and _4896_(_2465_, _2464_, encrypting);
    and _4897_(_2466_, _2465_, _0781_);
    and _4898_(_2467_, _0799_, cipher_key[92]);
    or _4899_(_2468_, _2467_, _2466_);
    and _4900_(_2469_, _2468_, _0794_);
    or _4901_(_0611_, _2469_, _2463_);
    and _4902_(_2470_, _0792_, round_key[93]);
    and _4903_(_2471_, _0779_, round_key[85]);
    and _4904_(_2472_, _2471_, encrypting);
    and _4905_(_2473_, _2472_, _0781_);
    and _4906_(_2474_, _0799_, cipher_key[93]);
    or _4907_(_2475_, _2474_, _2473_);
    and _4908_(_2476_, _2475_, _0794_);
    or _4909_(_0612_, _2476_, _2470_);
    and _4910_(_2477_, _0792_, round_key[94]);
    and _4911_(_2478_, _0779_, round_key[86]);
    and _4912_(_2479_, _2478_, encrypting);
    and _4913_(_2480_, _2479_, _0781_);
    and _4914_(_2481_, _0799_, cipher_key[94]);
    or _4915_(_2482_, _2481_, _2480_);
    and _4916_(_2483_, _2482_, _0794_);
    or _4917_(_0613_, _2483_, _2477_);
    and _4918_(_2484_, _0792_, round_key[95]);
    and _4919_(_2485_, _0779_, round_key[87]);
    and _4920_(_2486_, _2485_, encrypting);
    and _4921_(_2487_, _2486_, _0781_);
    and _4922_(_2488_, _0799_, cipher_key[95]);
    or _4923_(_2489_, _2488_, _2487_);
    and _4924_(_2490_, _2489_, _0794_);
    or _4925_(_0614_, _2490_, _2484_);
    and _4926_(_2491_, _0792_, round_key[96]);
    and _4927_(_2492_, _0779_, round_key[88]);
    and _4928_(_2493_, _2492_, encrypting);
    and _4929_(_2494_, _2493_, _0781_);
    and _4930_(_2495_, _0799_, cipher_key[96]);
    or _4931_(_2496_, _2495_, _2494_);
    and _4932_(_2497_, _2496_, _0794_);
    or _4933_(_0615_, _2497_, _2491_);
    and _4934_(_2498_, _0792_, round_key[97]);
    and _4935_(_2499_, _0779_, round_key[89]);
    and _4936_(_2500_, _2499_, encrypting);
    and _4937_(_2501_, _2500_, _0781_);
    and _4938_(_2502_, _0799_, cipher_key[97]);
    or _4939_(_2503_, _2502_, _2501_);
    and _4940_(_2504_, _2503_, _0794_);
    or _4941_(_0616_, _2504_, _2498_);
    and _4942_(_2505_, _0792_, round_key[98]);
    and _4943_(_2506_, _0779_, round_key[90]);
    and _4944_(_2507_, _2506_, encrypting);
    and _4945_(_2508_, _2507_, _0781_);
    and _4946_(_2509_, _0799_, cipher_key[98]);
    or _4947_(_2510_, _2509_, _2508_);
    and _4948_(_2511_, _2510_, _0794_);
    or _4949_(_0617_, _2511_, _2505_);
    and _4950_(_2512_, _0792_, round_key[99]);
    and _4951_(_2513_, _0779_, round_key[91]);
    and _4952_(_2514_, _2513_, encrypting);
    and _4953_(_2515_, _2514_, _0781_);
    and _4954_(_2516_, _0799_, cipher_key[99]);
    or _4955_(_2517_, _2516_, _2515_);
    and _4956_(_2518_, _2517_, _0794_);
    or _4957_(_0618_, _2518_, _2512_);
    and _4958_(_2519_, _0792_, round_key[100]);
    and _4959_(_2520_, _0779_, round_key[92]);
    and _4960_(_2521_, _2520_, encrypting);
    and _4961_(_2522_, _2521_, _0781_);
    and _4962_(_2523_, _0799_, cipher_key[100]);
    or _4963_(_2524_, _2523_, _2522_);
    and _4964_(_2525_, _2524_, _0794_);
    or _4965_(_0619_, _2525_, _2519_);
    and _4966_(_2526_, _0792_, round_key[101]);
    and _4967_(_2527_, _0779_, round_key[93]);
    and _4968_(_2528_, _2527_, encrypting);
    and _4969_(_2529_, _2528_, _0781_);
    and _4970_(_2530_, _0799_, cipher_key[101]);
    or _4971_(_2531_, _2530_, _2529_);
    and _4972_(_2532_, _2531_, _0794_);
    or _4973_(_0620_, _2532_, _2526_);
    and _4974_(_2533_, _0792_, round_key[102]);
    and _4975_(_2534_, _0779_, round_key[94]);
    and _4976_(_2535_, _2534_, encrypting);
    and _4977_(_2536_, _2535_, _0781_);
    and _4978_(_2537_, _0799_, cipher_key[102]);
    or _4979_(_2538_, _2537_, _2536_);
    and _4980_(_2539_, _2538_, _0794_);
    or _4981_(_0621_, _2539_, _2533_);
    and _4982_(_2540_, _0792_, round_key[103]);
    and _4983_(_2541_, _0779_, round_key[95]);
    and _4984_(_2542_, _2541_, encrypting);
    and _4985_(_2543_, _2542_, _0781_);
    and _4986_(_2544_, _0799_, cipher_key[103]);
    or _4987_(_2545_, _2544_, _2543_);
    and _4988_(_2546_, _2545_, _0794_);
    or _4989_(_0622_, _2546_, _2540_);
    and _4990_(_2547_, _0792_, round_key[104]);
    and _4991_(_2548_, _0779_, round_key[96]);
    and _4992_(_2549_, _2548_, encrypting);
    and _4993_(_2550_, _2549_, _0781_);
    and _4994_(_2551_, _0799_, cipher_key[104]);
    or _4995_(_2552_, _2551_, _2550_);
    and _4996_(_2553_, _2552_, _0794_);
    or _4997_(_0623_, _2553_, _2547_);
    and _4998_(_2554_, _0792_, round_key[105]);
    and _4999_(_2555_, _0779_, round_key[97]);
    and _5000_(_2556_, _2555_, encrypting);
    and _5001_(_2557_, _2556_, _0781_);
    and _5002_(_2558_, _0799_, cipher_key[105]);
    or _5003_(_2559_, _2558_, _2557_);
    and _5004_(_2560_, _2559_, _0794_);
    or _5005_(_0624_, _2560_, _2554_);
    and _5006_(_2561_, _0792_, round_key[106]);
    and _5007_(_2562_, _0779_, round_key[98]);
    and _5008_(_2563_, _2562_, encrypting);
    and _5009_(_2564_, _2563_, _0781_);
    and _5010_(_2565_, _0799_, cipher_key[106]);
    or _5011_(_2566_, _2565_, _2564_);
    and _5012_(_2567_, _2566_, _0794_);
    or _5013_(_0625_, _2567_, _2561_);
    and _5014_(_2568_, _0792_, round_key[107]);
    and _5015_(_2569_, _0779_, round_key[99]);
    and _5016_(_2570_, _2569_, encrypting);
    and _5017_(_2571_, _2570_, _0781_);
    and _5018_(_2572_, _0799_, cipher_key[107]);
    or _5019_(_2573_, _2572_, _2571_);
    and _5020_(_2574_, _2573_, _0794_);
    or _5021_(_0626_, _2574_, _2568_);
    and _5022_(_2575_, _0792_, round_key[108]);
    and _5023_(_2576_, _0779_, round_key[100]);
    and _5024_(_2577_, _2576_, encrypting);
    and _5025_(_2578_, _2577_, _0781_);
    and _5026_(_2579_, _0799_, cipher_key[108]);
    or _5027_(_2580_, _2579_, _2578_);
    and _5028_(_2581_, _2580_, _0794_);
    or _5029_(_0627_, _2581_, _2575_);
    and _5030_(_2582_, _0792_, round_key[109]);
    and _5031_(_2583_, _0779_, round_key[101]);
    and _5032_(_2584_, _2583_, encrypting);
    and _5033_(_2585_, _2584_, _0781_);
    and _5034_(_2586_, _0799_, cipher_key[109]);
    or _5035_(_2587_, _2586_, _2585_);
    and _5036_(_2588_, _2587_, _0794_);
    or _5037_(_0628_, _2588_, _2582_);
    and _5038_(_2589_, _0792_, round_key[110]);
    and _5039_(_2590_, _0779_, round_key[102]);
    and _5040_(_2591_, _2590_, encrypting);
    and _5041_(_2592_, _2591_, _0781_);
    and _5042_(_2593_, _0799_, cipher_key[110]);
    or _5043_(_2594_, _2593_, _2592_);
    and _5044_(_2595_, _2594_, _0794_);
    or _5045_(_0629_, _2595_, _2589_);
    and _5046_(_2596_, _0792_, round_key[111]);
    and _5047_(_2597_, _0779_, round_key[103]);
    and _5048_(_2598_, _2597_, encrypting);
    and _5049_(_2599_, _2598_, _0781_);
    and _5050_(_2600_, _0799_, cipher_key[111]);
    or _5051_(_2601_, _2600_, _2599_);
    and _5052_(_2602_, _2601_, _0794_);
    or _5053_(_0630_, _2602_, _2596_);
    and _5054_(_2603_, _0792_, round_key[112]);
    and _5055_(_2604_, _0779_, round_key[104]);
    and _5056_(_2605_, _2604_, encrypting);
    and _5057_(_2606_, _2605_, _0781_);
    and _5058_(_2607_, _0799_, cipher_key[112]);
    or _5059_(_2608_, _2607_, _2606_);
    and _5060_(_2609_, _2608_, _0794_);
    or _5061_(_0631_, _2609_, _2603_);
    and _5062_(_2610_, _0792_, round_key[113]);
    and _5063_(_2611_, _0779_, round_key[105]);
    and _5064_(_2612_, _2611_, encrypting);
    and _5065_(_2613_, _2612_, _0781_);
    and _5066_(_2614_, _0799_, cipher_key[113]);
    or _5067_(_2615_, _2614_, _2613_);
    and _5068_(_2616_, _2615_, _0794_);
    or _5069_(_0632_, _2616_, _2610_);
    and _5070_(_2617_, _0792_, round_key[114]);
    and _5071_(_2618_, _0779_, round_key[106]);
    and _5072_(_2619_, _2618_, encrypting);
    and _5073_(_2620_, _2619_, _0781_);
    and _5074_(_2621_, _0799_, cipher_key[114]);
    or _5075_(_2622_, _2621_, _2620_);
    and _5076_(_2623_, _2622_, _0794_);
    or _5077_(_0633_, _2623_, _2617_);
    and _5078_(_2624_, _0792_, round_key[115]);
    and _5079_(_2625_, _0779_, round_key[107]);
    and _5080_(_2626_, _2625_, encrypting);
    and _5081_(_2627_, _2626_, _0781_);
    and _5082_(_2628_, _0799_, cipher_key[115]);
    or _5083_(_2629_, _2628_, _2627_);
    and _5084_(_2630_, _2629_, _0794_);
    or _5085_(_0634_, _2630_, _2624_);
    and _5086_(_2631_, _0792_, round_key[116]);
    and _5087_(_2632_, _0779_, round_key[108]);
    and _5088_(_2633_, _2632_, encrypting);
    and _5089_(_2634_, _2633_, _0781_);
    and _5090_(_2635_, _0799_, cipher_key[116]);
    or _5091_(_2636_, _2635_, _2634_);
    and _5092_(_2637_, _2636_, _0794_);
    or _5093_(_0635_, _2637_, _2631_);
    and _5094_(_2638_, _0792_, round_key[117]);
    and _5095_(_2639_, _0779_, round_key[109]);
    and _5096_(_2640_, _2639_, encrypting);
    and _5097_(_2641_, _2640_, _0781_);
    and _5098_(_2642_, _0799_, cipher_key[117]);
    or _5099_(_2643_, _2642_, _2641_);
    and _5100_(_2644_, _2643_, _0794_);
    or _5101_(_0636_, _2644_, _2638_);
    and _5102_(_2645_, _0792_, round_key[118]);
    and _5103_(_2646_, _0779_, round_key[110]);
    and _5104_(_2647_, _2646_, encrypting);
    and _5105_(_2648_, _2647_, _0781_);
    and _5106_(_2649_, _0799_, cipher_key[118]);
    or _5107_(_2650_, _2649_, _2648_);
    and _5108_(_2651_, _2650_, _0794_);
    or _5109_(_0637_, _2651_, _2645_);
    and _5110_(_2652_, _0792_, round_key[119]);
    and _5111_(_2653_, _0779_, round_key[111]);
    and _5112_(_2654_, _2653_, encrypting);
    and _5113_(_2655_, _2654_, _0781_);
    and _5114_(_2656_, _0799_, cipher_key[119]);
    or _5115_(_2657_, _2656_, _2655_);
    and _5116_(_2658_, _2657_, _0794_);
    or _5117_(_0638_, _2658_, _2652_);
    and _5118_(_2659_, _0792_, round_key[120]);
    and _5119_(_2660_, _0779_, round_key[112]);
    and _5120_(_2661_, _2660_, encrypting);
    and _5121_(_2662_, _2661_, _0781_);
    and _5122_(_2663_, _0799_, cipher_key[120]);
    or _5123_(_2664_, _2663_, _2662_);
    and _5124_(_2665_, _2664_, _0794_);
    or _5125_(_0639_, _2665_, _2659_);
    and _5126_(_2666_, _0792_, round_key[121]);
    and _5127_(_2667_, _0779_, round_key[113]);
    and _5128_(_2668_, _2667_, encrypting);
    and _5129_(_2669_, _2668_, _0781_);
    and _5130_(_2670_, _0799_, cipher_key[121]);
    or _5131_(_2671_, _2670_, _2669_);
    and _5132_(_2672_, _2671_, _0794_);
    or _5133_(_0640_, _2672_, _2666_);
    and _5134_(_2673_, _0792_, round_key[122]);
    and _5135_(_2674_, _0779_, round_key[114]);
    and _5136_(_2675_, _2674_, encrypting);
    and _5137_(_2676_, _2675_, _0781_);
    and _5138_(_2677_, _0799_, cipher_key[122]);
    or _5139_(_2678_, _2677_, _2676_);
    and _5140_(_2679_, _2678_, _0794_);
    or _5141_(_0641_, _2679_, _2673_);
    and _5142_(_2680_, _0792_, round_key[123]);
    and _5143_(_2681_, _0779_, round_key[115]);
    and _5144_(_2682_, _2681_, encrypting);
    and _5145_(_2683_, _2682_, _0781_);
    and _5146_(_2684_, _0799_, cipher_key[123]);
    or _5147_(_2685_, _2684_, _2683_);
    and _5148_(_2686_, _2685_, _0794_);
    or _5149_(_0642_, _2686_, _2680_);
    and _5150_(_2687_, _0792_, round_key[124]);
    and _5151_(_2688_, _0779_, round_key[116]);
    and _5152_(_2689_, _2688_, encrypting);
    and _5153_(_2690_, _2689_, _0781_);
    and _5154_(_2691_, _0799_, cipher_key[124]);
    or _5155_(_2692_, _2691_, _2690_);
    and _5156_(_2693_, _2692_, _0794_);
    or _5157_(_0643_, _2693_, _2687_);
    and _5158_(_2694_, _0792_, round_key[125]);
    and _5159_(_2695_, _0779_, round_key[117]);
    and _5160_(_2696_, _2695_, encrypting);
    and _5161_(_2697_, _2696_, _0781_);
    and _5162_(_2698_, _0799_, cipher_key[125]);
    or _5163_(_2699_, _2698_, _2697_);
    and _5164_(_2700_, _2699_, _0794_);
    or _5165_(_0644_, _2700_, _2694_);
    and _5166_(_2701_, _0792_, round_key[126]);
    and _5167_(_2702_, _0779_, round_key[118]);
    and _5168_(_2703_, _2702_, encrypting);
    and _5169_(_2704_, _2703_, _0781_);
    and _5170_(_2705_, _0799_, cipher_key[126]);
    or _5171_(_2706_, _2705_, _2704_);
    and _5172_(_2707_, _2706_, _0794_);
    or _5173_(_0645_, _2707_, _2701_);
    and _5174_(_2708_, _0792_, round_key[127]);
    and _5175_(_2709_, _0779_, round_key[119]);
    and _5176_(_2710_, _2709_, encrypting);
    and _5177_(_2711_, _2710_, _0781_);
    and _5178_(_2712_, _0799_, cipher_key[127]);
    or _5179_(_2713_, _2712_, _2711_);
    and _5180_(_2714_, _2713_, _0794_);
    or _5181_(_0646_, _2714_, _2708_);
    and _5182_(_2715_, _0792_, round_counter[0]);
    nor _5183_(_2716_, _0785_, round_counter[0]);
    and _5184_(_2717_, _2716_, encrypting);
    and _5185_(_2718_, _2717_, _0781_);
    and _5186_(_2719_, _2718_, _0794_);
    or _5187_(_0647_, _2719_, _2715_);
    and _5188_(_2720_, _0792_, round_counter[1]);
    xor _5189_(_2721_, round_counter[1], round_counter[0]);
    and _5190_(_2722_, _2721_, encrypting);
    and _5191_(_2723_, _2722_, _0781_);
    and _5192_(_2724_, _2723_, _0794_);
    or _5193_(_0648_, _2724_, _2720_);
    and _5194_(_2725_, _0792_, round_counter[2]);
    xor _5195_(_2726_, _0778_, round_counter[2]);
    and _5196_(_2727_, _2726_, encrypting);
    and _5197_(_2728_, _2727_, _0781_);
    and _5198_(_2729_, _2728_, _0794_);
    or _5199_(_0649_, _2729_, _2725_);
    and _5200_(_2730_, _0788_, ciphertext[0]);
    and _5201_(_2731_, _0787_, state[0]);
    or _5202_(_0650_, _2731_, _2730_);
    and _5203_(_2732_, _0788_, ciphertext[1]);
    and _5204_(_2733_, _0787_, state[1]);
    or _5205_(_0651_, _2733_, _2732_);
    and _5206_(_2734_, _0788_, ciphertext[2]);
    and _5207_(_2735_, _0787_, state[2]);
    or _5208_(_0652_, _2735_, _2734_);
    and _5209_(_2736_, _0788_, ciphertext[3]);
    and _5210_(_2737_, _0787_, state[3]);
    or _5211_(_0653_, _2737_, _2736_);
    and _5212_(_2738_, _0788_, ciphertext[4]);
    and _5213_(_2739_, _0787_, state[4]);
    or _5214_(_0654_, _2739_, _2738_);
    and _5215_(_2740_, _0788_, ciphertext[5]);
    and _5216_(_2741_, _0787_, state[5]);
    or _5217_(_0655_, _2741_, _2740_);
    and _5218_(_2742_, _0788_, ciphertext[6]);
    and _5219_(_2743_, _0787_, state[6]);
    or _5220_(_0656_, _2743_, _2742_);
    and _5221_(_2744_, _0788_, ciphertext[7]);
    and _5222_(_2745_, _0787_, state[7]);
    or _5223_(_0657_, _2745_, _2744_);
    and _5224_(_2746_, _0788_, ciphertext[8]);
    and _5225_(_2747_, _0787_, state[8]);
    or _5226_(_0658_, _2747_, _2746_);
    and _5227_(_2748_, _0788_, ciphertext[9]);
    and _5228_(_2749_, _0787_, state[9]);
    or _5229_(_0659_, _2749_, _2748_);
    and _5230_(_2750_, _0788_, ciphertext[10]);
    and _5231_(_2751_, _0787_, state[10]);
    or _5232_(_0660_, _2751_, _2750_);
    and _5233_(_2752_, _0788_, ciphertext[11]);
    and _5234_(_2753_, _0787_, state[11]);
    or _5235_(_0661_, _2753_, _2752_);
    and _5236_(_2754_, _0788_, ciphertext[12]);
    and _5237_(_2755_, _0787_, state[12]);
    or _5238_(_0662_, _2755_, _2754_);
    and _5239_(_2756_, _0788_, ciphertext[13]);
    and _5240_(_2757_, _0787_, state[13]);
    or _5241_(_0663_, _2757_, _2756_);
    and _5242_(_2758_, _0788_, ciphertext[14]);
    and _5243_(_2759_, _0787_, state[14]);
    or _5244_(_0664_, _2759_, _2758_);
    and _5245_(_2760_, _0788_, ciphertext[15]);
    and _5246_(_2761_, _0787_, state[15]);
    or _5247_(_0665_, _2761_, _2760_);
    and _5248_(_2762_, _0788_, ciphertext[16]);
    and _5249_(_2763_, _0787_, state[16]);
    or _5250_(_0666_, _2763_, _2762_);
    and _5251_(_2764_, _0788_, ciphertext[17]);
    and _5252_(_2765_, _0787_, state[17]);
    or _5253_(_0667_, _2765_, _2764_);
    and _5254_(_2766_, _0788_, ciphertext[18]);
    and _5255_(_2767_, _0787_, state[18]);
    or _5256_(_0668_, _2767_, _2766_);
    and _5257_(_2768_, _0788_, ciphertext[19]);
    and _5258_(_2769_, _0787_, state[19]);
    or _5259_(_0669_, _2769_, _2768_);
    and _5260_(_2770_, _0788_, ciphertext[20]);
    and _5261_(_2771_, _0787_, state[20]);
    or _5262_(_0670_, _2771_, _2770_);
    and _5263_(_2772_, _0788_, ciphertext[21]);
    and _5264_(_2773_, _0787_, state[21]);
    or _5265_(_0671_, _2773_, _2772_);
    and _5266_(_2774_, _0788_, ciphertext[22]);
    and _5267_(_2775_, _0787_, state[22]);
    or _5268_(_0672_, _2775_, _2774_);
    and _5269_(_2776_, _0788_, ciphertext[23]);
    and _5270_(_2777_, _0787_, state[23]);
    or _5271_(_0673_, _2777_, _2776_);
    and _5272_(_2778_, _0788_, ciphertext[24]);
    and _5273_(_2779_, _0787_, state[24]);
    or _5274_(_0674_, _2779_, _2778_);
    and _5275_(_2780_, _0788_, ciphertext[25]);
    and _5276_(_2781_, _0787_, state[25]);
    or _5277_(_0675_, _2781_, _2780_);
    and _5278_(_2782_, _0788_, ciphertext[26]);
    and _5279_(_2783_, _0787_, state[26]);
    or _5280_(_0676_, _2783_, _2782_);
    and _5281_(_2784_, _0788_, ciphertext[27]);
    and _5282_(_2785_, _0787_, state[27]);
    or _5283_(_0677_, _2785_, _2784_);
    and _5284_(_2786_, _0788_, ciphertext[28]);
    and _5285_(_2787_, _0787_, state[28]);
    or _5286_(_0678_, _2787_, _2786_);
    and _5287_(_2788_, _0788_, ciphertext[29]);
    and _5288_(_2789_, _0787_, state[29]);
    or _5289_(_0679_, _2789_, _2788_);
    and _5290_(_2790_, _0788_, ciphertext[30]);
    and _5291_(_2791_, _0787_, state[30]);
    or _5292_(_0680_, _2791_, _2790_);
    and _5293_(_2792_, _0788_, ciphertext[31]);
    and _5294_(_2793_, _0787_, state[31]);
    or _5295_(_0681_, _2793_, _2792_);
    and _5296_(_2794_, _0788_, ciphertext[32]);
    and _5297_(_2795_, _0787_, state[32]);
    or _5298_(_0682_, _2795_, _2794_);
    and _5299_(_2796_, _0788_, ciphertext[33]);
    and _5300_(_2797_, _0787_, state[33]);
    or _5301_(_0683_, _2797_, _2796_);
    and _5302_(_2798_, _0788_, ciphertext[34]);
    and _5303_(_2799_, _0787_, state[34]);
    or _5304_(_0684_, _2799_, _2798_);
    and _5305_(_2800_, _0788_, ciphertext[35]);
    and _5306_(_2801_, _0787_, state[35]);
    or _5307_(_0685_, _2801_, _2800_);
    and _5308_(_2802_, _0788_, ciphertext[36]);
    and _5309_(_2803_, _0787_, state[36]);
    or _5310_(_0686_, _2803_, _2802_);
    and _5311_(_2804_, _0788_, ciphertext[37]);
    and _5312_(_2805_, _0787_, state[37]);
    or _5313_(_0687_, _2805_, _2804_);
    and _5314_(_2806_, _0788_, ciphertext[38]);
    and _5315_(_2807_, _0787_, state[38]);
    or _5316_(_0688_, _2807_, _2806_);
    and _5317_(_2808_, _0788_, ciphertext[39]);
    and _5318_(_2809_, _0787_, state[39]);
    or _5319_(_0689_, _2809_, _2808_);
    and _5320_(_2810_, _0788_, ciphertext[40]);
    and _5321_(_2811_, _0787_, state[40]);
    or _5322_(_0690_, _2811_, _2810_);
    and _5323_(_2812_, _0788_, ciphertext[41]);
    and _5324_(_2813_, _0787_, state[41]);
    or _5325_(_0691_, _2813_, _2812_);
    and _5326_(_2814_, _0788_, ciphertext[42]);
    and _5327_(_2815_, _0787_, state[42]);
    or _5328_(_0692_, _2815_, _2814_);
    and _5329_(_2816_, _0788_, ciphertext[43]);
    and _5330_(_2817_, _0787_, state[43]);
    or _5331_(_0693_, _2817_, _2816_);
    and _5332_(_2818_, _0788_, ciphertext[44]);
    and _5333_(_2819_, _0787_, state[44]);
    or _5334_(_0694_, _2819_, _2818_);
    and _5335_(_2820_, _0788_, ciphertext[45]);
    and _5336_(_2821_, _0787_, state[45]);
    or _5337_(_0695_, _2821_, _2820_);
    and _5338_(_2822_, _0788_, ciphertext[46]);
    and _5339_(_2823_, _0787_, state[46]);
    or _5340_(_0696_, _2823_, _2822_);
    and _5341_(_2824_, _0788_, ciphertext[47]);
    and _5342_(_2825_, _0787_, state[47]);
    or _5343_(_0697_, _2825_, _2824_);
    and _5344_(_2826_, _0788_, ciphertext[48]);
    and _5345_(_2827_, _0787_, state[48]);
    or _5346_(_0698_, _2827_, _2826_);
    and _5347_(_2828_, _0788_, ciphertext[49]);
    and _5348_(_2829_, _0787_, state[49]);
    or _5349_(_0699_, _2829_, _2828_);
    and _5350_(_2830_, _0788_, ciphertext[50]);
    and _5351_(_2831_, _0787_, state[50]);
    or _5352_(_0700_, _2831_, _2830_);
    and _5353_(_2832_, _0788_, ciphertext[51]);
    and _5354_(_2833_, _0787_, state[51]);
    or _5355_(_0701_, _2833_, _2832_);
    and _5356_(_2834_, _0788_, ciphertext[52]);
    and _5357_(_2835_, _0787_, state[52]);
    or _5358_(_0702_, _2835_, _2834_);
    and _5359_(_2836_, _0788_, ciphertext[53]);
    and _5360_(_2837_, _0787_, state[53]);
    or _5361_(_0703_, _2837_, _2836_);
    and _5362_(_2838_, _0788_, ciphertext[54]);
    and _5363_(_2839_, _0787_, state[54]);
    or _5364_(_0704_, _2839_, _2838_);
    and _5365_(_2840_, _0788_, ciphertext[55]);
    and _5366_(_2841_, _0787_, state[55]);
    or _5367_(_0705_, _2841_, _2840_);
    and _5368_(_2842_, _0788_, ciphertext[56]);
    and _5369_(_2843_, _0787_, state[56]);
    or _5370_(_0706_, _2843_, _2842_);
    and _5371_(_2844_, _0788_, ciphertext[57]);
    and _5372_(_2845_, _0787_, state[57]);
    or _5373_(_0707_, _2845_, _2844_);
    and _5374_(_2846_, _0788_, ciphertext[58]);
    and _5375_(_2847_, _0787_, state[58]);
    or _5376_(_0708_, _2847_, _2846_);
    and _5377_(_2848_, _0788_, ciphertext[59]);
    and _5378_(_2849_, _0787_, state[59]);
    or _5379_(_0709_, _2849_, _2848_);
    and _5380_(_2850_, _0788_, ciphertext[60]);
    and _5381_(_2851_, _0787_, state[60]);
    or _5382_(_0710_, _2851_, _2850_);
    and _5383_(_2852_, _0788_, ciphertext[61]);
    and _5384_(_2853_, _0787_, state[61]);
    or _5385_(_0711_, _2853_, _2852_);
    and _5386_(_2854_, _0788_, ciphertext[62]);
    and _5387_(_2855_, _0787_, state[62]);
    or _5388_(_0712_, _2855_, _2854_);
    and _5389_(_2856_, _0788_, ciphertext[63]);
    and _5390_(_2857_, _0787_, state[63]);
    or _5391_(_0713_, _2857_, _2856_);
    and _5392_(_2858_, _0788_, ciphertext[64]);
    and _5393_(_2859_, _0787_, state[64]);
    or _5394_(_0714_, _2859_, _2858_);
    and _5395_(_2860_, _0788_, ciphertext[65]);
    and _5396_(_2861_, _0787_, state[65]);
    or _5397_(_0715_, _2861_, _2860_);
    and _5398_(_2862_, _0788_, ciphertext[66]);
    and _5399_(_2863_, _0787_, state[66]);
    or _5400_(_0716_, _2863_, _2862_);
    and _5401_(_2864_, _0788_, ciphertext[67]);
    and _5402_(_2865_, _0787_, state[67]);
    or _5403_(_0717_, _2865_, _2864_);
    and _5404_(_2866_, _0788_, ciphertext[68]);
    and _5405_(_2867_, _0787_, state[68]);
    or _5406_(_0718_, _2867_, _2866_);
    and _5407_(_2868_, _0788_, ciphertext[69]);
    and _5408_(_2869_, _0787_, state[69]);
    or _5409_(_0719_, _2869_, _2868_);
    and _5410_(_2870_, _0788_, ciphertext[70]);
    and _5411_(_2871_, _0787_, state[70]);
    or _5412_(_0720_, _2871_, _2870_);
    and _5413_(_2872_, _0788_, ciphertext[71]);
    and _5414_(_2873_, _0787_, state[71]);
    or _5415_(_0721_, _2873_, _2872_);
    and _5416_(_2874_, _0788_, ciphertext[72]);
    and _5417_(_2875_, _0787_, state[72]);
    or _5418_(_0722_, _2875_, _2874_);
    and _5419_(_2876_, _0788_, ciphertext[73]);
    and _5420_(_2877_, _0787_, state[73]);
    or _5421_(_0723_, _2877_, _2876_);
    and _5422_(_2878_, _0788_, ciphertext[74]);
    and _5423_(_2879_, _0787_, state[74]);
    or _5424_(_0724_, _2879_, _2878_);
    and _5425_(_2880_, _0788_, ciphertext[75]);
    and _5426_(_2881_, _0787_, state[75]);
    or _5427_(_0725_, _2881_, _2880_);
    and _5428_(_2882_, _0788_, ciphertext[76]);
    and _5429_(_2883_, _0787_, state[76]);
    or _5430_(_0726_, _2883_, _2882_);
    and _5431_(_2884_, _0788_, ciphertext[77]);
    and _5432_(_2885_, _0787_, state[77]);
    or _5433_(_0727_, _2885_, _2884_);
    and _5434_(_2886_, _0788_, ciphertext[78]);
    and _5435_(_2887_, _0787_, state[78]);
    or _5436_(_0728_, _2887_, _2886_);
    and _5437_(_2888_, _0788_, ciphertext[79]);
    and _5438_(_2889_, _0787_, state[79]);
    or _5439_(_0729_, _2889_, _2888_);
    and _5440_(_2890_, _0788_, ciphertext[80]);
    and _5441_(_2891_, _0787_, state[80]);
    or _5442_(_0730_, _2891_, _2890_);
    and _5443_(_2892_, _0788_, ciphertext[81]);
    and _5444_(_2893_, _0787_, state[81]);
    or _5445_(_0731_, _2893_, _2892_);
    and _5446_(_2894_, _0788_, ciphertext[82]);
    and _5447_(_2895_, _0787_, state[82]);
    or _5448_(_0732_, _2895_, _2894_);
    and _5449_(_2896_, _0788_, ciphertext[83]);
    and _5450_(_2897_, _0787_, state[83]);
    or _5451_(_0733_, _2897_, _2896_);
    and _5452_(_2898_, _0788_, ciphertext[84]);
    and _5453_(_2899_, _0787_, state[84]);
    or _5454_(_0734_, _2899_, _2898_);
    and _5455_(_2900_, _0788_, ciphertext[85]);
    and _5456_(_2901_, _0787_, state[85]);
    or _5457_(_0735_, _2901_, _2900_);
    and _5458_(_2902_, _0788_, ciphertext[86]);
    and _5459_(_2903_, _0787_, state[86]);
    or _5460_(_0736_, _2903_, _2902_);
    and _5461_(_2904_, _0788_, ciphertext[87]);
    and _5462_(_2905_, _0787_, state[87]);
    or _5463_(_0737_, _2905_, _2904_);
    and _5464_(_2906_, _0788_, ciphertext[88]);
    and _5465_(_2907_, _0787_, state[88]);
    or _5466_(_0738_, _2907_, _2906_);
    and _5467_(_2908_, _0788_, ciphertext[89]);
    and _5468_(_2909_, _0787_, state[89]);
    or _5469_(_0739_, _2909_, _2908_);
    and _5470_(_2910_, _0788_, ciphertext[90]);
    and _5471_(_2911_, _0787_, state[90]);
    or _5472_(_0740_, _2911_, _2910_);
    and _5473_(_2912_, _0788_, ciphertext[91]);
    and _5474_(_2913_, _0787_, state[91]);
    or _5475_(_0741_, _2913_, _2912_);
    and _5476_(_2914_, _0788_, ciphertext[92]);
    and _5477_(_2915_, _0787_, state[92]);
    or _5478_(_0742_, _2915_, _2914_);
    and _5479_(_2916_, _0788_, ciphertext[93]);
    and _5480_(_2917_, _0787_, state[93]);
    or _5481_(_0743_, _2917_, _2916_);
    and _5482_(_2918_, _0788_, ciphertext[94]);
    and _5483_(_2919_, _0787_, state[94]);
    or _5484_(_0744_, _2919_, _2918_);
    and _5485_(_2920_, _0788_, ciphertext[95]);
    and _5486_(_2921_, _0787_, state[95]);
    or _5487_(_0745_, _2921_, _2920_);
    and _5488_(_2922_, _0788_, ciphertext[96]);
    and _5489_(_2923_, _0787_, state[96]);
    or _5490_(_0746_, _2923_, _2922_);
    and _5491_(_2924_, _0788_, ciphertext[97]);
    and _5492_(_2925_, _0787_, state[97]);
    or _5493_(_0747_, _2925_, _2924_);
    and _5494_(_2926_, _0788_, ciphertext[98]);
    and _5495_(_2927_, _0787_, state[98]);
    or _5496_(_0748_, _2927_, _2926_);
    and _5497_(_2928_, _0788_, ciphertext[99]);
    and _5498_(_2929_, _0787_, state[99]);
    or _5499_(_0749_, _2929_, _2928_);
    and _5500_(_2930_, _0788_, ciphertext[100]);
    and _5501_(_2931_, _0787_, state[100]);
    or _5502_(_0750_, _2931_, _2930_);
    and _5503_(_2932_, _0788_, ciphertext[101]);
    and _5504_(_2933_, _0787_, state[101]);
    or _5505_(_0751_, _2933_, _2932_);
    and _5506_(_2934_, _0788_, ciphertext[102]);
    and _5507_(_2935_, _0787_, state[102]);
    or _5508_(_0752_, _2935_, _2934_);
    and _5509_(_2936_, _0788_, ciphertext[103]);
    and _5510_(_2937_, _0787_, state[103]);
    or _5511_(_0753_, _2937_, _2936_);
    and _5512_(_2938_, _0788_, ciphertext[104]);
    and _5513_(_2939_, _0787_, state[104]);
    or _5514_(_0754_, _2939_, _2938_);
    and _5515_(_2940_, _0788_, ciphertext[105]);
    and _5516_(_2941_, _0787_, state[105]);
    or _5517_(_0755_, _2941_, _2940_);
    and _5518_(_2942_, _0788_, ciphertext[106]);
    and _5519_(_2943_, _0787_, state[106]);
    or _5520_(_0756_, _2943_, _2942_);
    and _5521_(_2944_, _0788_, ciphertext[107]);
    and _5522_(_2945_, _0787_, state[107]);
    or _5523_(_0757_, _2945_, _2944_);
    and _5524_(_2946_, _0788_, ciphertext[108]);
    and _5525_(_2947_, _0787_, state[108]);
    or _5526_(_0758_, _2947_, _2946_);
    and _5527_(_2948_, _0788_, ciphertext[109]);
    and _5528_(_2949_, _0787_, state[109]);
    or _5529_(_0759_, _2949_, _2948_);
    and _5530_(_2950_, _0788_, ciphertext[110]);
    and _5531_(_2951_, _0787_, state[110]);
    or _5532_(_0760_, _2951_, _2950_);
    and _5533_(_2952_, _0788_, ciphertext[111]);
    and _5534_(_2953_, _0787_, state[111]);
    or _5535_(_0761_, _2953_, _2952_);
    and _5536_(_2954_, _0788_, ciphertext[112]);
    and _5537_(_2955_, _0787_, state[112]);
    or _5538_(_0762_, _2955_, _2954_);
    and _5539_(_2956_, _0788_, ciphertext[113]);
    and _5540_(_2957_, _0787_, state[113]);
    or _5541_(_0763_, _2957_, _2956_);
    and _5542_(_2958_, _0788_, ciphertext[114]);
    and _5543_(_2959_, _0787_, state[114]);
    or _5544_(_0764_, _2959_, _2958_);
    and _5545_(_2960_, _0788_, ciphertext[115]);
    and _5546_(_2961_, _0787_, state[115]);
    or _5547_(_0765_, _2961_, _2960_);
    and _5548_(_2962_, _0788_, ciphertext[116]);
    and _5549_(_2963_, _0787_, state[116]);
    or _5550_(_0766_, _2963_, _2962_);
    and _5551_(_2964_, _0788_, ciphertext[117]);
    and _5552_(_2965_, _0787_, state[117]);
    or _5553_(_0767_, _2965_, _2964_);
    and _5554_(_2966_, _0788_, ciphertext[118]);
    and _5555_(_2967_, _0787_, state[118]);
    or _5556_(_0768_, _2967_, _2966_);
    and _5557_(_2968_, _0788_, ciphertext[119]);
    and _5558_(_2969_, _0787_, state[119]);
    or _5559_(_0769_, _2969_, _2968_);
    and _5560_(_2970_, _0788_, ciphertext[120]);
    and _5561_(_2971_, _0787_, state[120]);
    or _5562_(_0770_, _2971_, _2970_);
    and _5563_(_2972_, _0788_, ciphertext[121]);
    and _5564_(_2973_, _0787_, state[121]);
    or _5565_(_0771_, _2973_, _2972_);
    and _5566_(_2974_, _0788_, ciphertext[122]);
    and _5567_(_2975_, _0787_, state[122]);
    or _5568_(_0772_, _2975_, _2974_);
    and _5569_(_2976_, _0788_, ciphertext[123]);
    and _5570_(_2977_, _0787_, state[123]);
    or _5571_(_0773_, _2977_, _2976_);
    and _5572_(_2978_, _0788_, ciphertext[124]);
    and _5573_(_2979_, _0787_, state[124]);
    or _5574_(_0774_, _2979_, _2978_);
    and _5575_(_2980_, _0788_, ciphertext[125]);
    and _5576_(_2981_, _0787_, state[125]);
    or _5577_(_0775_, _2981_, _2980_);
    and _5578_(_2982_, _0788_, ciphertext[126]);
    and _5579_(_2983_, _0787_, state[126]);
    or _5580_(_0776_, _2983_, _2982_);
    and _5581_(_2984_, _0788_, ciphertext[127]);
    and _5582_(_2985_, _0787_, state[127]);
    or _5583_(_0777_, _2985_, _2984_);
    and _5584_(_2986_, _0779_, encrypting);
    or _5585_(_0000_, _2986_, _0799_);
    not _5586_(_0002_, rst);
    not _5587_(_0003_, rst);
    not _5588_(_0004_, rst);
    not _5589_(_0005_, rst);
    not _5590_(_0006_, rst);
    not _5591_(_0007_, rst);
    not _5592_(_0008_, rst);
    not _5593_(_0009_, rst);
    not _5594_(_0010_, rst);
    not _5595_(_0011_, rst);
    not _5596_(_0012_, rst);
    not _5597_(_0013_, rst);
    not _5598_(_0014_, rst);
    not _5599_(_0015_, rst);
    not _5600_(_0016_, rst);
    not _5601_(_0017_, rst);
    not _5602_(_0018_, rst);
    not _5603_(_0019_, rst);
    not _5604_(_0020_, rst);
    not _5605_(_0021_, rst);
    not _5606_(_0022_, rst);
    not _5607_(_0023_, rst);
    not _5608_(_0024_, rst);
    not _5609_(_0025_, rst);
    not _5610_(_0026_, rst);
    not _5611_(_0027_, rst);
    not _5612_(_0028_, rst);
    not _5613_(_0029_, rst);
    not _5614_(_0030_, rst);
    not _5615_(_0031_, rst);
    not _5616_(_0032_, rst);
    not _5617_(_0033_, rst);
    not _5618_(_0034_, rst);
    not _5619_(_0035_, rst);
    not _5620_(_0036_, rst);
    not _5621_(_0037_, rst);
    not _5622_(_0038_, rst);
    not _5623_(_0039_, rst);
    not _5624_(_0040_, rst);
    not _5625_(_0041_, rst);
    not _5626_(_0042_, rst);
    not _5627_(_0043_, rst);
    not _5628_(_0044_, rst);
    not _5629_(_0045_, rst);
    not _5630_(_0046_, rst);
    not _5631_(_0047_, rst);
    not _5632_(_0048_, rst);
    not _5633_(_0049_, rst);
    not _5634_(_0050_, rst);
    not _5635_(_0051_, rst);
    not _5636_(_0052_, rst);
    not _5637_(_0053_, rst);
    not _5638_(_0054_, rst);
    not _5639_(_0055_, rst);
    not _5640_(_0056_, rst);
    not _5641_(_0057_, rst);
    not _5642_(_0058_, rst);
    not _5643_(_0059_, rst);
    not _5644_(_0060_, rst);
    not _5645_(_0061_, rst);
    not _5646_(_0062_, rst);
    not _5647_(_0063_, rst);
    not _5648_(_0064_, rst);
    not _5649_(_0065_, rst);
    not _5650_(_0066_, rst);
    not _5651_(_0067_, rst);
    not _5652_(_0068_, rst);
    not _5653_(_0069_, rst);
    not _5654_(_0070_, rst);
    not _5655_(_0071_, rst);
    not _5656_(_0072_, rst);
    not _5657_(_0073_, rst);
    not _5658_(_0074_, rst);
    not _5659_(_0075_, rst);
    not _5660_(_0076_, rst);
    not _5661_(_0077_, rst);
    not _5662_(_0078_, rst);
    not _5663_(_0079_, rst);
    not _5664_(_0080_, rst);
    not _5665_(_0081_, rst);
    not _5666_(_0082_, rst);
    not _5667_(_0083_, rst);
    not _5668_(_0084_, rst);
    not _5669_(_0085_, rst);
    not _5670_(_0086_, rst);
    not _5671_(_0087_, rst);
    not _5672_(_0088_, rst);
    not _5673_(_0089_, rst);
    not _5674_(_0090_, rst);
    not _5675_(_0091_, rst);
    not _5676_(_0092_, rst);
    not _5677_(_0093_, rst);
    not _5678_(_0094_, rst);
    not _5679_(_0095_, rst);
    not _5680_(_0096_, rst);
    not _5681_(_0097_, rst);
    not _5682_(_0098_, rst);
    not _5683_(_0099_, rst);
    not _5684_(_0100_, rst);
    not _5685_(_0101_, rst);
    not _5686_(_0102_, rst);
    not _5687_(_0103_, rst);
    not _5688_(_0104_, rst);
    not _5689_(_0105_, rst);
    not _5690_(_0106_, rst);
    not _5691_(_0107_, rst);
    not _5692_(_0108_, rst);
    not _5693_(_0109_, rst);
    not _5694_(_0110_, rst);
    not _5695_(_0111_, rst);
    not _5696_(_0112_, rst);
    not _5697_(_0113_, rst);
    not _5698_(_0114_, rst);
    not _5699_(_0115_, rst);
    not _5700_(_0116_, rst);
    not _5701_(_0117_, rst);
    not _5702_(_0118_, rst);
    not _5703_(_0119_, rst);
    not _5704_(_0120_, rst);
    not _5705_(_0121_, rst);
    not _5706_(_0122_, rst);
    not _5707_(_0123_, rst);
    not _5708_(_0124_, rst);
    not _5709_(_0125_, rst);
    not _5710_(_0126_, rst);
    not _5711_(_0127_, rst);
    not _5712_(_0128_, rst);
    not _5713_(_0129_, rst);
    not _5714_(_0130_, rst);
    not _5715_(_0131_, rst);
    not _5716_(_0132_, rst);
    not _5717_(_0133_, rst);
    not _5718_(_0134_, rst);
    not _5719_(_0135_, rst);
    not _5720_(_0136_, rst);
    not _5721_(_0137_, rst);
    not _5722_(_0138_, rst);
    not _5723_(_0139_, rst);
    not _5724_(_0140_, rst);
    not _5725_(_0141_, rst);
    not _5726_(_0142_, rst);
    not _5727_(_0143_, rst);
    not _5728_(_0144_, rst);
    not _5729_(_0145_, rst);
    not _5730_(_0146_, rst);
    not _5731_(_0147_, rst);
    not _5732_(_0148_, rst);
    not _5733_(_0149_, rst);
    not _5734_(_0150_, rst);
    not _5735_(_0151_, rst);
    not _5736_(_0152_, rst);
    not _5737_(_0153_, rst);
    not _5738_(_0154_, rst);
    not _5739_(_0155_, rst);
    not _5740_(_0156_, rst);
    not _5741_(_0157_, rst);
    not _5742_(_0158_, rst);
    not _5743_(_0159_, rst);
    not _5744_(_0160_, rst);
    not _5745_(_0161_, rst);
    not _5746_(_0162_, rst);
    not _5747_(_0163_, rst);
    not _5748_(_0164_, rst);
    not _5749_(_0165_, rst);
    not _5750_(_0166_, rst);
    not _5751_(_0167_, rst);
    not _5752_(_0168_, rst);
    not _5753_(_0169_, rst);
    not _5754_(_0170_, rst);
    not _5755_(_0171_, rst);
    not _5756_(_0172_, rst);
    not _5757_(_0173_, rst);
    not _5758_(_0174_, rst);
    not _5759_(_0175_, rst);
    not _5760_(_0176_, rst);
    not _5761_(_0177_, rst);
    not _5762_(_0178_, rst);
    not _5763_(_0179_, rst);
    not _5764_(_0180_, rst);
    not _5765_(_0181_, rst);
    not _5766_(_0182_, rst);
    not _5767_(_0183_, rst);
    not _5768_(_0184_, rst);
    not _5769_(_0185_, rst);
    not _5770_(_0186_, rst);
    not _5771_(_0187_, rst);
    not _5772_(_0188_, rst);
    not _5773_(_0189_, rst);
    not _5774_(_0190_, rst);
    not _5775_(_0191_, rst);
    not _5776_(_0192_, rst);
    not _5777_(_0193_, rst);
    not _5778_(_0194_, rst);
    not _5779_(_0195_, rst);
    not _5780_(_0196_, rst);
    not _5781_(_0197_, rst);
    not _5782_(_0198_, rst);
    not _5783_(_0199_, rst);
    not _5784_(_0200_, rst);
    not _5785_(_0201_, rst);
    not _5786_(_0202_, rst);
    not _5787_(_0203_, rst);
    not _5788_(_0204_, rst);
    not _5789_(_0205_, rst);
    not _5790_(_0206_, rst);
    not _5791_(_0207_, rst);
    not _5792_(_0208_, rst);
    not _5793_(_0209_, rst);
    not _5794_(_0210_, rst);
    not _5795_(_0211_, rst);
    not _5796_(_0212_, rst);
    not _5797_(_0213_, rst);
    not _5798_(_0214_, rst);
    not _5799_(_0215_, rst);
    not _5800_(_0216_, rst);
    not _5801_(_0217_, rst);
    not _5802_(_0218_, rst);
    not _5803_(_0219_, rst);
    not _5804_(_0220_, rst);
    not _5805_(_0221_, rst);
    not _5806_(_0222_, rst);
    not _5807_(_0223_, rst);
    not _5808_(_0224_, rst);
    not _5809_(_0225_, rst);
    not _5810_(_0226_, rst);
    not _5811_(_0227_, rst);
    not _5812_(_0228_, rst);
    not _5813_(_0229_, rst);
    not _5814_(_0230_, rst);
    not _5815_(_0231_, rst);
    not _5816_(_0232_, rst);
    not _5817_(_0233_, rst);
    not _5818_(_0234_, rst);
    not _5819_(_0235_, rst);
    not _5820_(_0236_, rst);
    not _5821_(_0237_, rst);
    not _5822_(_0238_, rst);
    not _5823_(_0239_, rst);
    not _5824_(_0240_, rst);
    not _5825_(_0241_, rst);
    not _5826_(_0242_, rst);
    not _5827_(_0243_, rst);
    not _5828_(_0244_, rst);
    not _5829_(_0245_, rst);
    not _5830_(_0246_, rst);
    not _5831_(_0247_, rst);
    not _5832_(_0248_, rst);
    not _5833_(_0249_, rst);
    not _5834_(_0250_, rst);
    not _5835_(_0251_, rst);
    not _5836_(_0252_, rst);
    not _5837_(_0253_, rst);
    not _5838_(_0254_, rst);
    not _5839_(_0255_, rst);
    not _5840_(_0256_, rst);
    not _5841_(_0257_, rst);
    not _5842_(_0258_, rst);
    not _5843_(_0259_, rst);
    not _5844_(_0260_, rst);
    not _5845_(_0261_, rst);
    not _5846_(_0262_, rst);
    not _5847_(_0263_, rst);
    not _5848_(_0264_, rst);
    not _5849_(_0265_, rst);
    not _5850_(_0266_, rst);
    not _5851_(_0267_, rst);
    not _5852_(_0268_, rst);
    not _5853_(_0269_, rst);
    not _5854_(_0270_, rst);
    not _5855_(_0271_, rst);
    not _5856_(_0272_, rst);
    not _5857_(_0273_, rst);
    not _5858_(_0274_, rst);
    not _5859_(_0275_, rst);
    not _5860_(_0276_, rst);
    not _5861_(_0277_, rst);
    not _5862_(_0278_, rst);
    not _5863_(_0279_, rst);
    not _5864_(_0280_, rst);
    not _5865_(_0281_, rst);
    not _5866_(_0282_, rst);
    not _5867_(_0283_, rst);
    not _5868_(_0284_, rst);
    not _5869_(_0285_, rst);
    not _5870_(_0286_, rst);
    not _5871_(_0287_, rst);
    not _5872_(_0288_, rst);
    not _5873_(_0289_, rst);
    not _5874_(_0290_, rst);
    not _5875_(_0291_, rst);
    not _5876_(_0292_, rst);
    not _5877_(_0293_, rst);
    not _5878_(_0294_, rst);
    not _5879_(_0295_, rst);
    not _5880_(_0296_, rst);
    not _5881_(_0297_, rst);
    not _5882_(_0298_, rst);
    not _5883_(_0299_, rst);
    not _5884_(_0300_, rst);
    not _5885_(_0301_, rst);
    not _5886_(_0302_, rst);
    not _5887_(_0303_, rst);
    not _5888_(_0304_, rst);
    not _5889_(_0305_, rst);
    not _5890_(_0306_, rst);
    not _5891_(_0307_, rst);
    not _5892_(_0308_, rst);
    not _5893_(_0309_, rst);
    not _5894_(_0310_, rst);
    not _5895_(_0311_, rst);
    not _5896_(_0312_, rst);
    not _5897_(_0313_, rst);
    not _5898_(_0314_, rst);
    not _5899_(_0315_, rst);
    not _5900_(_0316_, rst);
    not _5901_(_0317_, rst);
    not _5902_(_0318_, rst);
    not _5903_(_0319_, rst);
    not _5904_(_0320_, rst);
    not _5905_(_0321_, rst);
    not _5906_(_0322_, rst);
    not _5907_(_0323_, rst);
    not _5908_(_0324_, rst);
    not _5909_(_0325_, rst);
    not _5910_(_0326_, rst);
    not _5911_(_0327_, rst);
    not _5912_(_0328_, rst);
    not _5913_(_0329_, rst);
    not _5914_(_0330_, rst);
    not _5915_(_0331_, rst);
    not _5916_(_0332_, rst);
    not _5917_(_0333_, rst);
    not _5918_(_0334_, rst);
    not _5919_(_0335_, rst);
    not _5920_(_0336_, rst);
    not _5921_(_0337_, rst);
    not _5922_(_0338_, rst);
    not _5923_(_0339_, rst);
    not _5924_(_0340_, rst);
    not _5925_(_0341_, rst);
    not _5926_(_0342_, rst);
    not _5927_(_0343_, rst);
    not _5928_(_0344_, rst);
    not _5929_(_0345_, rst);
    not _5930_(_0346_, rst);
    not _5931_(_0347_, rst);
    not _5932_(_0348_, rst);
    not _5933_(_0349_, rst);
    not _5934_(_0350_, rst);
    not _5935_(_0351_, rst);
    not _5936_(_0352_, rst);
    not _5937_(_0353_, rst);
    not _5938_(_0354_, rst);
    not _5939_(_0355_, rst);
    not _5940_(_0356_, rst);
    not _5941_(_0357_, rst);
    not _5942_(_0358_, rst);
    not _5943_(_0359_, rst);
    not _5944_(_0360_, rst);
    not _5945_(_0361_, rst);
    not _5946_(_0362_, rst);
    not _5947_(_0363_, rst);
    not _5948_(_0364_, rst);
    not _5949_(_0365_, rst);
    not _5950_(_0366_, rst);
    not _5951_(_0367_, rst);
    not _5952_(_0368_, rst);
    not _5953_(_0369_, rst);
    not _5954_(_0370_, rst);
    not _5955_(_0371_, rst);
    not _5956_(_0372_, rst);
    not _5957_(_0373_, rst);
    not _5958_(_0374_, rst);
    not _5959_(_0375_, rst);
    not _5960_(_0376_, rst);
    not _5961_(_0377_, rst);
    not _5962_(_0378_, rst);
    not _5963_(_0379_, rst);
    not _5964_(_0380_, rst);
    not _5965_(_0381_, rst);
    not _5966_(_0382_, rst);
    not _5967_(_0383_, rst);
    not _5968_(_0384_, rst);
    not _5969_(_0385_, rst);
    not _5970_(_0386_, rst);
    not _5971_(_0387_, rst);
    not _5972_(_0388_, rst);
    not _5973_(_0389_, rst);
    dff _5974_(.RN(_0001_), .SN(1'b1), .CK(clk), .D(_0390_), .Q(encrypt_done));
    dff _5975_(.RN(_0002_), .SN(1'b1), .CK(clk), .D(_0391_), .Q(state[0]));
    dff _5976_(.RN(_0003_), .SN(1'b1), .CK(clk), .D(_0392_), .Q(state[1]));
    dff _5977_(.RN(_0004_), .SN(1'b1), .CK(clk), .D(_0393_), .Q(state[2]));
    dff _5978_(.RN(_0005_), .SN(1'b1), .CK(clk), .D(_0394_), .Q(state[3]));
    dff _5979_(.RN(_0006_), .SN(1'b1), .CK(clk), .D(_0395_), .Q(state[4]));
    dff _5980_(.RN(_0007_), .SN(1'b1), .CK(clk), .D(_0396_), .Q(state[5]));
    dff _5981_(.RN(_0008_), .SN(1'b1), .CK(clk), .D(_0397_), .Q(state[6]));
    dff _5982_(.RN(_0009_), .SN(1'b1), .CK(clk), .D(_0398_), .Q(state[7]));
    dff _5983_(.RN(_0010_), .SN(1'b1), .CK(clk), .D(_0399_), .Q(state[8]));
    dff _5984_(.RN(_0011_), .SN(1'b1), .CK(clk), .D(_0400_), .Q(state[9]));
    dff _5985_(.RN(_0012_), .SN(1'b1), .CK(clk), .D(_0401_), .Q(state[10]));
    dff _5986_(.RN(_0013_), .SN(1'b1), .CK(clk), .D(_0402_), .Q(state[11]));
    dff _5987_(.RN(_0014_), .SN(1'b1), .CK(clk), .D(_0403_), .Q(state[12]));
    dff _5988_(.RN(_0015_), .SN(1'b1), .CK(clk), .D(_0404_), .Q(state[13]));
    dff _5989_(.RN(_0016_), .SN(1'b1), .CK(clk), .D(_0405_), .Q(state[14]));
    dff _5990_(.RN(_0017_), .SN(1'b1), .CK(clk), .D(_0406_), .Q(state[15]));
    dff _5991_(.RN(_0018_), .SN(1'b1), .CK(clk), .D(_0407_), .Q(state[16]));
    dff _5992_(.RN(_0019_), .SN(1'b1), .CK(clk), .D(_0408_), .Q(state[17]));
    dff _5993_(.RN(_0020_), .SN(1'b1), .CK(clk), .D(_0409_), .Q(state[18]));
    dff _5994_(.RN(_0021_), .SN(1'b1), .CK(clk), .D(_0410_), .Q(state[19]));
    dff _5995_(.RN(_0022_), .SN(1'b1), .CK(clk), .D(_0411_), .Q(state[20]));
    dff _5996_(.RN(_0023_), .SN(1'b1), .CK(clk), .D(_0412_), .Q(state[21]));
    dff _5997_(.RN(_0024_), .SN(1'b1), .CK(clk), .D(_0413_), .Q(state[22]));
    dff _5998_(.RN(_0025_), .SN(1'b1), .CK(clk), .D(_0414_), .Q(state[23]));
    dff _5999_(.RN(_0026_), .SN(1'b1), .CK(clk), .D(_0415_), .Q(state[24]));
    dff _6000_(.RN(_0027_), .SN(1'b1), .CK(clk), .D(_0416_), .Q(state[25]));
    dff _6001_(.RN(_0028_), .SN(1'b1), .CK(clk), .D(_0417_), .Q(state[26]));
    dff _6002_(.RN(_0029_), .SN(1'b1), .CK(clk), .D(_0418_), .Q(state[27]));
    dff _6003_(.RN(_0030_), .SN(1'b1), .CK(clk), .D(_0419_), .Q(state[28]));
    dff _6004_(.RN(_0031_), .SN(1'b1), .CK(clk), .D(_0420_), .Q(state[29]));
    dff _6005_(.RN(_0032_), .SN(1'b1), .CK(clk), .D(_0421_), .Q(state[30]));
    dff _6006_(.RN(_0033_), .SN(1'b1), .CK(clk), .D(_0422_), .Q(state[31]));
    dff _6007_(.RN(_0034_), .SN(1'b1), .CK(clk), .D(_0423_), .Q(state[32]));
    dff _6008_(.RN(_0035_), .SN(1'b1), .CK(clk), .D(_0424_), .Q(state[33]));
    dff _6009_(.RN(_0036_), .SN(1'b1), .CK(clk), .D(_0425_), .Q(state[34]));
    dff _6010_(.RN(_0037_), .SN(1'b1), .CK(clk), .D(_0426_), .Q(state[35]));
    dff _6011_(.RN(_0038_), .SN(1'b1), .CK(clk), .D(_0427_), .Q(state[36]));
    dff _6012_(.RN(_0039_), .SN(1'b1), .CK(clk), .D(_0428_), .Q(state[37]));
    dff _6013_(.RN(_0040_), .SN(1'b1), .CK(clk), .D(_0429_), .Q(state[38]));
    dff _6014_(.RN(_0041_), .SN(1'b1), .CK(clk), .D(_0430_), .Q(state[39]));
    dff _6015_(.RN(_0042_), .SN(1'b1), .CK(clk), .D(_0431_), .Q(state[40]));
    dff _6016_(.RN(_0043_), .SN(1'b1), .CK(clk), .D(_0432_), .Q(state[41]));
    dff _6017_(.RN(_0044_), .SN(1'b1), .CK(clk), .D(_0433_), .Q(state[42]));
    dff _6018_(.RN(_0045_), .SN(1'b1), .CK(clk), .D(_0434_), .Q(state[43]));
    dff _6019_(.RN(_0046_), .SN(1'b1), .CK(clk), .D(_0435_), .Q(state[44]));
    dff _6020_(.RN(_0047_), .SN(1'b1), .CK(clk), .D(_0436_), .Q(state[45]));
    dff _6021_(.RN(_0048_), .SN(1'b1), .CK(clk), .D(_0437_), .Q(state[46]));
    dff _6022_(.RN(_0049_), .SN(1'b1), .CK(clk), .D(_0438_), .Q(state[47]));
    dff _6023_(.RN(_0050_), .SN(1'b1), .CK(clk), .D(_0439_), .Q(state[48]));
    dff _6024_(.RN(_0051_), .SN(1'b1), .CK(clk), .D(_0440_), .Q(state[49]));
    dff _6025_(.RN(_0052_), .SN(1'b1), .CK(clk), .D(_0441_), .Q(state[50]));
    dff _6026_(.RN(_0053_), .SN(1'b1), .CK(clk), .D(_0442_), .Q(state[51]));
    dff _6027_(.RN(_0054_), .SN(1'b1), .CK(clk), .D(_0443_), .Q(state[52]));
    dff _6028_(.RN(_0055_), .SN(1'b1), .CK(clk), .D(_0444_), .Q(state[53]));
    dff _6029_(.RN(_0056_), .SN(1'b1), .CK(clk), .D(_0445_), .Q(state[54]));
    dff _6030_(.RN(_0057_), .SN(1'b1), .CK(clk), .D(_0446_), .Q(state[55]));
    dff _6031_(.RN(_0058_), .SN(1'b1), .CK(clk), .D(_0447_), .Q(state[56]));
    dff _6032_(.RN(_0059_), .SN(1'b1), .CK(clk), .D(_0448_), .Q(state[57]));
    dff _6033_(.RN(_0060_), .SN(1'b1), .CK(clk), .D(_0449_), .Q(state[58]));
    dff _6034_(.RN(_0061_), .SN(1'b1), .CK(clk), .D(_0450_), .Q(state[59]));
    dff _6035_(.RN(_0062_), .SN(1'b1), .CK(clk), .D(_0451_), .Q(state[60]));
    dff _6036_(.RN(_0063_), .SN(1'b1), .CK(clk), .D(_0452_), .Q(state[61]));
    dff _6037_(.RN(_0064_), .SN(1'b1), .CK(clk), .D(_0453_), .Q(state[62]));
    dff _6038_(.RN(_0065_), .SN(1'b1), .CK(clk), .D(_0454_), .Q(state[63]));
    dff _6039_(.RN(_0066_), .SN(1'b1), .CK(clk), .D(_0455_), .Q(state[64]));
    dff _6040_(.RN(_0067_), .SN(1'b1), .CK(clk), .D(_0456_), .Q(state[65]));
    dff _6041_(.RN(_0068_), .SN(1'b1), .CK(clk), .D(_0457_), .Q(state[66]));
    dff _6042_(.RN(_0069_), .SN(1'b1), .CK(clk), .D(_0458_), .Q(state[67]));
    dff _6043_(.RN(_0070_), .SN(1'b1), .CK(clk), .D(_0459_), .Q(state[68]));
    dff _6044_(.RN(_0071_), .SN(1'b1), .CK(clk), .D(_0460_), .Q(state[69]));
    dff _6045_(.RN(_0072_), .SN(1'b1), .CK(clk), .D(_0461_), .Q(state[70]));
    dff _6046_(.RN(_0073_), .SN(1'b1), .CK(clk), .D(_0462_), .Q(state[71]));
    dff _6047_(.RN(_0074_), .SN(1'b1), .CK(clk), .D(_0463_), .Q(state[72]));
    dff _6048_(.RN(_0075_), .SN(1'b1), .CK(clk), .D(_0464_), .Q(state[73]));
    dff _6049_(.RN(_0076_), .SN(1'b1), .CK(clk), .D(_0465_), .Q(state[74]));
    dff _6050_(.RN(_0077_), .SN(1'b1), .CK(clk), .D(_0466_), .Q(state[75]));
    dff _6051_(.RN(_0078_), .SN(1'b1), .CK(clk), .D(_0467_), .Q(state[76]));
    dff _6052_(.RN(_0079_), .SN(1'b1), .CK(clk), .D(_0468_), .Q(state[77]));
    dff _6053_(.RN(_0080_), .SN(1'b1), .CK(clk), .D(_0469_), .Q(state[78]));
    dff _6054_(.RN(_0081_), .SN(1'b1), .CK(clk), .D(_0470_), .Q(state[79]));
    dff _6055_(.RN(_0082_), .SN(1'b1), .CK(clk), .D(_0471_), .Q(state[80]));
    dff _6056_(.RN(_0083_), .SN(1'b1), .CK(clk), .D(_0472_), .Q(state[81]));
    dff _6057_(.RN(_0084_), .SN(1'b1), .CK(clk), .D(_0473_), .Q(state[82]));
    dff _6058_(.RN(_0085_), .SN(1'b1), .CK(clk), .D(_0474_), .Q(state[83]));
    dff _6059_(.RN(_0086_), .SN(1'b1), .CK(clk), .D(_0475_), .Q(state[84]));
    dff _6060_(.RN(_0087_), .SN(1'b1), .CK(clk), .D(_0476_), .Q(state[85]));
    dff _6061_(.RN(_0088_), .SN(1'b1), .CK(clk), .D(_0477_), .Q(state[86]));
    dff _6062_(.RN(_0089_), .SN(1'b1), .CK(clk), .D(_0478_), .Q(state[87]));
    dff _6063_(.RN(_0090_), .SN(1'b1), .CK(clk), .D(_0479_), .Q(state[88]));
    dff _6064_(.RN(_0091_), .SN(1'b1), .CK(clk), .D(_0480_), .Q(state[89]));
    dff _6065_(.RN(_0092_), .SN(1'b1), .CK(clk), .D(_0481_), .Q(state[90]));
    dff _6066_(.RN(_0093_), .SN(1'b1), .CK(clk), .D(_0482_), .Q(state[91]));
    dff _6067_(.RN(_0094_), .SN(1'b1), .CK(clk), .D(_0483_), .Q(state[92]));
    dff _6068_(.RN(_0095_), .SN(1'b1), .CK(clk), .D(_0484_), .Q(state[93]));
    dff _6069_(.RN(_0096_), .SN(1'b1), .CK(clk), .D(_0485_), .Q(state[94]));
    dff _6070_(.RN(_0097_), .SN(1'b1), .CK(clk), .D(_0486_), .Q(state[95]));
    dff _6071_(.RN(_0098_), .SN(1'b1), .CK(clk), .D(_0487_), .Q(state[96]));
    dff _6072_(.RN(_0099_), .SN(1'b1), .CK(clk), .D(_0488_), .Q(state[97]));
    dff _6073_(.RN(_0100_), .SN(1'b1), .CK(clk), .D(_0489_), .Q(state[98]));
    dff _6074_(.RN(_0101_), .SN(1'b1), .CK(clk), .D(_0490_), .Q(state[99]));
    dff _6075_(.RN(_0102_), .SN(1'b1), .CK(clk), .D(_0491_), .Q(state[100]));
    dff _6076_(.RN(_0103_), .SN(1'b1), .CK(clk), .D(_0492_), .Q(state[101]));
    dff _6077_(.RN(_0104_), .SN(1'b1), .CK(clk), .D(_0493_), .Q(state[102]));
    dff _6078_(.RN(_0105_), .SN(1'b1), .CK(clk), .D(_0494_), .Q(state[103]));
    dff _6079_(.RN(_0106_), .SN(1'b1), .CK(clk), .D(_0495_), .Q(state[104]));
    dff _6080_(.RN(_0107_), .SN(1'b1), .CK(clk), .D(_0496_), .Q(state[105]));
    dff _6081_(.RN(_0108_), .SN(1'b1), .CK(clk), .D(_0497_), .Q(state[106]));
    dff _6082_(.RN(_0109_), .SN(1'b1), .CK(clk), .D(_0498_), .Q(state[107]));
    dff _6083_(.RN(_0110_), .SN(1'b1), .CK(clk), .D(_0499_), .Q(state[108]));
    dff _6084_(.RN(_0111_), .SN(1'b1), .CK(clk), .D(_0500_), .Q(state[109]));
    dff _6085_(.RN(_0112_), .SN(1'b1), .CK(clk), .D(_0501_), .Q(state[110]));
    dff _6086_(.RN(_0113_), .SN(1'b1), .CK(clk), .D(_0502_), .Q(state[111]));
    dff _6087_(.RN(_0114_), .SN(1'b1), .CK(clk), .D(_0503_), .Q(state[112]));
    dff _6088_(.RN(_0115_), .SN(1'b1), .CK(clk), .D(_0504_), .Q(state[113]));
    dff _6089_(.RN(_0116_), .SN(1'b1), .CK(clk), .D(_0505_), .Q(state[114]));
    dff _6090_(.RN(_0117_), .SN(1'b1), .CK(clk), .D(_0506_), .Q(state[115]));
    dff _6091_(.RN(_0118_), .SN(1'b1), .CK(clk), .D(_0507_), .Q(state[116]));
    dff _6092_(.RN(_0119_), .SN(1'b1), .CK(clk), .D(_0508_), .Q(state[117]));
    dff _6093_(.RN(_0120_), .SN(1'b1), .CK(clk), .D(_0509_), .Q(state[118]));
    dff _6094_(.RN(_0121_), .SN(1'b1), .CK(clk), .D(_0510_), .Q(state[119]));
    dff _6095_(.RN(_0122_), .SN(1'b1), .CK(clk), .D(_0511_), .Q(state[120]));
    dff _6096_(.RN(_0123_), .SN(1'b1), .CK(clk), .D(_0512_), .Q(state[121]));
    dff _6097_(.RN(_0124_), .SN(1'b1), .CK(clk), .D(_0513_), .Q(state[122]));
    dff _6098_(.RN(_0125_), .SN(1'b1), .CK(clk), .D(_0514_), .Q(state[123]));
    dff _6099_(.RN(_0126_), .SN(1'b1), .CK(clk), .D(_0515_), .Q(state[124]));
    dff _6100_(.RN(_0127_), .SN(1'b1), .CK(clk), .D(_0516_), .Q(state[125]));
    dff _6101_(.RN(_0128_), .SN(1'b1), .CK(clk), .D(_0517_), .Q(state[126]));
    dff _6102_(.RN(_0129_), .SN(1'b1), .CK(clk), .D(_0518_), .Q(state[127]));
    dff _6103_(.RN(_0130_), .SN(1'b1), .CK(clk), .D(_0519_), .Q(round_key[0]));
    dff _6104_(.RN(_0131_), .SN(1'b1), .CK(clk), .D(_0520_), .Q(round_key[1]));
    dff _6105_(.RN(_0132_), .SN(1'b1), .CK(clk), .D(_0521_), .Q(round_key[2]));
    dff _6106_(.RN(_0133_), .SN(1'b1), .CK(clk), .D(_0522_), .Q(round_key[3]));
    dff _6107_(.RN(_0134_), .SN(1'b1), .CK(clk), .D(_0523_), .Q(round_key[4]));
    dff _6108_(.RN(_0135_), .SN(1'b1), .CK(clk), .D(_0524_), .Q(round_key[5]));
    dff _6109_(.RN(_0136_), .SN(1'b1), .CK(clk), .D(_0525_), .Q(round_key[6]));
    dff _6110_(.RN(_0137_), .SN(1'b1), .CK(clk), .D(_0526_), .Q(round_key[7]));
    dff _6111_(.RN(_0138_), .SN(1'b1), .CK(clk), .D(_0527_), .Q(round_key[8]));
    dff _6112_(.RN(_0139_), .SN(1'b1), .CK(clk), .D(_0528_), .Q(round_key[9]));
    dff _6113_(.RN(_0140_), .SN(1'b1), .CK(clk), .D(_0529_), .Q(round_key[10]));
    dff _6114_(.RN(_0141_), .SN(1'b1), .CK(clk), .D(_0530_), .Q(round_key[11]));
    dff _6115_(.RN(_0142_), .SN(1'b1), .CK(clk), .D(_0531_), .Q(round_key[12]));
    dff _6116_(.RN(_0143_), .SN(1'b1), .CK(clk), .D(_0532_), .Q(round_key[13]));
    dff _6117_(.RN(_0144_), .SN(1'b1), .CK(clk), .D(_0533_), .Q(round_key[14]));
    dff _6118_(.RN(_0145_), .SN(1'b1), .CK(clk), .D(_0534_), .Q(round_key[15]));
    dff _6119_(.RN(_0146_), .SN(1'b1), .CK(clk), .D(_0535_), .Q(round_key[16]));
    dff _6120_(.RN(_0147_), .SN(1'b1), .CK(clk), .D(_0536_), .Q(round_key[17]));
    dff _6121_(.RN(_0148_), .SN(1'b1), .CK(clk), .D(_0537_), .Q(round_key[18]));
    dff _6122_(.RN(_0149_), .SN(1'b1), .CK(clk), .D(_0538_), .Q(round_key[19]));
    dff _6123_(.RN(_0150_), .SN(1'b1), .CK(clk), .D(_0539_), .Q(round_key[20]));
    dff _6124_(.RN(_0151_), .SN(1'b1), .CK(clk), .D(_0540_), .Q(round_key[21]));
    dff _6125_(.RN(_0152_), .SN(1'b1), .CK(clk), .D(_0541_), .Q(round_key[22]));
    dff _6126_(.RN(_0153_), .SN(1'b1), .CK(clk), .D(_0542_), .Q(round_key[23]));
    dff _6127_(.RN(_0154_), .SN(1'b1), .CK(clk), .D(_0543_), .Q(round_key[24]));
    dff _6128_(.RN(_0155_), .SN(1'b1), .CK(clk), .D(_0544_), .Q(round_key[25]));
    dff _6129_(.RN(_0156_), .SN(1'b1), .CK(clk), .D(_0545_), .Q(round_key[26]));
    dff _6130_(.RN(_0157_), .SN(1'b1), .CK(clk), .D(_0546_), .Q(round_key[27]));
    dff _6131_(.RN(_0158_), .SN(1'b1), .CK(clk), .D(_0547_), .Q(round_key[28]));
    dff _6132_(.RN(_0159_), .SN(1'b1), .CK(clk), .D(_0548_), .Q(round_key[29]));
    dff _6133_(.RN(_0160_), .SN(1'b1), .CK(clk), .D(_0549_), .Q(round_key[30]));
    dff _6134_(.RN(_0161_), .SN(1'b1), .CK(clk), .D(_0550_), .Q(round_key[31]));
    dff _6135_(.RN(_0162_), .SN(1'b1), .CK(clk), .D(_0551_), .Q(round_key[32]));
    dff _6136_(.RN(_0163_), .SN(1'b1), .CK(clk), .D(_0552_), .Q(round_key[33]));
    dff _6137_(.RN(_0164_), .SN(1'b1), .CK(clk), .D(_0553_), .Q(round_key[34]));
    dff _6138_(.RN(_0165_), .SN(1'b1), .CK(clk), .D(_0554_), .Q(round_key[35]));
    dff _6139_(.RN(_0166_), .SN(1'b1), .CK(clk), .D(_0555_), .Q(round_key[36]));
    dff _6140_(.RN(_0167_), .SN(1'b1), .CK(clk), .D(_0556_), .Q(round_key[37]));
    dff _6141_(.RN(_0168_), .SN(1'b1), .CK(clk), .D(_0557_), .Q(round_key[38]));
    dff _6142_(.RN(_0169_), .SN(1'b1), .CK(clk), .D(_0558_), .Q(round_key[39]));
    dff _6143_(.RN(_0170_), .SN(1'b1), .CK(clk), .D(_0559_), .Q(round_key[40]));
    dff _6144_(.RN(_0171_), .SN(1'b1), .CK(clk), .D(_0560_), .Q(round_key[41]));
    dff _6145_(.RN(_0172_), .SN(1'b1), .CK(clk), .D(_0561_), .Q(round_key[42]));
    dff _6146_(.RN(_0173_), .SN(1'b1), .CK(clk), .D(_0562_), .Q(round_key[43]));
    dff _6147_(.RN(_0174_), .SN(1'b1), .CK(clk), .D(_0563_), .Q(round_key[44]));
    dff _6148_(.RN(_0175_), .SN(1'b1), .CK(clk), .D(_0564_), .Q(round_key[45]));
    dff _6149_(.RN(_0176_), .SN(1'b1), .CK(clk), .D(_0565_), .Q(round_key[46]));
    dff _6150_(.RN(_0177_), .SN(1'b1), .CK(clk), .D(_0566_), .Q(round_key[47]));
    dff _6151_(.RN(_0178_), .SN(1'b1), .CK(clk), .D(_0567_), .Q(round_key[48]));
    dff _6152_(.RN(_0179_), .SN(1'b1), .CK(clk), .D(_0568_), .Q(round_key[49]));
    dff _6153_(.RN(_0180_), .SN(1'b1), .CK(clk), .D(_0569_), .Q(round_key[50]));
    dff _6154_(.RN(_0181_), .SN(1'b1), .CK(clk), .D(_0570_), .Q(round_key[51]));
    dff _6155_(.RN(_0182_), .SN(1'b1), .CK(clk), .D(_0571_), .Q(round_key[52]));
    dff _6156_(.RN(_0183_), .SN(1'b1), .CK(clk), .D(_0572_), .Q(round_key[53]));
    dff _6157_(.RN(_0184_), .SN(1'b1), .CK(clk), .D(_0573_), .Q(round_key[54]));
    dff _6158_(.RN(_0185_), .SN(1'b1), .CK(clk), .D(_0574_), .Q(round_key[55]));
    dff _6159_(.RN(_0186_), .SN(1'b1), .CK(clk), .D(_0575_), .Q(round_key[56]));
    dff _6160_(.RN(_0187_), .SN(1'b1), .CK(clk), .D(_0576_), .Q(round_key[57]));
    dff _6161_(.RN(_0188_), .SN(1'b1), .CK(clk), .D(_0577_), .Q(round_key[58]));
    dff _6162_(.RN(_0189_), .SN(1'b1), .CK(clk), .D(_0578_), .Q(round_key[59]));
    dff _6163_(.RN(_0190_), .SN(1'b1), .CK(clk), .D(_0579_), .Q(round_key[60]));
    dff _6164_(.RN(_0191_), .SN(1'b1), .CK(clk), .D(_0580_), .Q(round_key[61]));
    dff _6165_(.RN(_0192_), .SN(1'b1), .CK(clk), .D(_0581_), .Q(round_key[62]));
    dff _6166_(.RN(_0193_), .SN(1'b1), .CK(clk), .D(_0582_), .Q(round_key[63]));
    dff _6167_(.RN(_0194_), .SN(1'b1), .CK(clk), .D(_0583_), .Q(round_key[64]));
    dff _6168_(.RN(_0195_), .SN(1'b1), .CK(clk), .D(_0584_), .Q(round_key[65]));
    dff _6169_(.RN(_0196_), .SN(1'b1), .CK(clk), .D(_0585_), .Q(round_key[66]));
    dff _6170_(.RN(_0197_), .SN(1'b1), .CK(clk), .D(_0586_), .Q(round_key[67]));
    dff _6171_(.RN(_0198_), .SN(1'b1), .CK(clk), .D(_0587_), .Q(round_key[68]));
    dff _6172_(.RN(_0199_), .SN(1'b1), .CK(clk), .D(_0588_), .Q(round_key[69]));
    dff _6173_(.RN(_0200_), .SN(1'b1), .CK(clk), .D(_0589_), .Q(round_key[70]));
    dff _6174_(.RN(_0201_), .SN(1'b1), .CK(clk), .D(_0590_), .Q(round_key[71]));
    dff _6175_(.RN(_0202_), .SN(1'b1), .CK(clk), .D(_0591_), .Q(round_key[72]));
    dff _6176_(.RN(_0203_), .SN(1'b1), .CK(clk), .D(_0592_), .Q(round_key[73]));
    dff _6177_(.RN(_0204_), .SN(1'b1), .CK(clk), .D(_0593_), .Q(round_key[74]));
    dff _6178_(.RN(_0205_), .SN(1'b1), .CK(clk), .D(_0594_), .Q(round_key[75]));
    dff _6179_(.RN(_0206_), .SN(1'b1), .CK(clk), .D(_0595_), .Q(round_key[76]));
    dff _6180_(.RN(_0207_), .SN(1'b1), .CK(clk), .D(_0596_), .Q(round_key[77]));
    dff _6181_(.RN(_0208_), .SN(1'b1), .CK(clk), .D(_0597_), .Q(round_key[78]));
    dff _6182_(.RN(_0209_), .SN(1'b1), .CK(clk), .D(_0598_), .Q(round_key[79]));
    dff _6183_(.RN(_0210_), .SN(1'b1), .CK(clk), .D(_0599_), .Q(round_key[80]));
    dff _6184_(.RN(_0211_), .SN(1'b1), .CK(clk), .D(_0600_), .Q(round_key[81]));
    dff _6185_(.RN(_0212_), .SN(1'b1), .CK(clk), .D(_0601_), .Q(round_key[82]));
    dff _6186_(.RN(_0213_), .SN(1'b1), .CK(clk), .D(_0602_), .Q(round_key[83]));
    dff _6187_(.RN(_0214_), .SN(1'b1), .CK(clk), .D(_0603_), .Q(round_key[84]));
    dff _6188_(.RN(_0215_), .SN(1'b1), .CK(clk), .D(_0604_), .Q(round_key[85]));
    dff _6189_(.RN(_0216_), .SN(1'b1), .CK(clk), .D(_0605_), .Q(round_key[86]));
    dff _6190_(.RN(_0217_), .SN(1'b1), .CK(clk), .D(_0606_), .Q(round_key[87]));
    dff _6191_(.RN(_0218_), .SN(1'b1), .CK(clk), .D(_0607_), .Q(round_key[88]));
    dff _6192_(.RN(_0219_), .SN(1'b1), .CK(clk), .D(_0608_), .Q(round_key[89]));
    dff _6193_(.RN(_0220_), .SN(1'b1), .CK(clk), .D(_0609_), .Q(round_key[90]));
    dff _6194_(.RN(_0221_), .SN(1'b1), .CK(clk), .D(_0610_), .Q(round_key[91]));
    dff _6195_(.RN(_0222_), .SN(1'b1), .CK(clk), .D(_0611_), .Q(round_key[92]));
    dff _6196_(.RN(_0223_), .SN(1'b1), .CK(clk), .D(_0612_), .Q(round_key[93]));
    dff _6197_(.RN(_0224_), .SN(1'b1), .CK(clk), .D(_0613_), .Q(round_key[94]));
    dff _6198_(.RN(_0225_), .SN(1'b1), .CK(clk), .D(_0614_), .Q(round_key[95]));
    dff _6199_(.RN(_0226_), .SN(1'b1), .CK(clk), .D(_0615_), .Q(round_key[96]));
    dff _6200_(.RN(_0227_), .SN(1'b1), .CK(clk), .D(_0616_), .Q(round_key[97]));
    dff _6201_(.RN(_0228_), .SN(1'b1), .CK(clk), .D(_0617_), .Q(round_key[98]));
    dff _6202_(.RN(_0229_), .SN(1'b1), .CK(clk), .D(_0618_), .Q(round_key[99]));
    dff _6203_(.RN(_0230_), .SN(1'b1), .CK(clk), .D(_0619_), .Q(round_key[100]));
    dff _6204_(.RN(_0231_), .SN(1'b1), .CK(clk), .D(_0620_), .Q(round_key[101]));
    dff _6205_(.RN(_0232_), .SN(1'b1), .CK(clk), .D(_0621_), .Q(round_key[102]));
    dff _6206_(.RN(_0233_), .SN(1'b1), .CK(clk), .D(_0622_), .Q(round_key[103]));
    dff _6207_(.RN(_0234_), .SN(1'b1), .CK(clk), .D(_0623_), .Q(round_key[104]));
    dff _6208_(.RN(_0235_), .SN(1'b1), .CK(clk), .D(_0624_), .Q(round_key[105]));
    dff _6209_(.RN(_0236_), .SN(1'b1), .CK(clk), .D(_0625_), .Q(round_key[106]));
    dff _6210_(.RN(_0237_), .SN(1'b1), .CK(clk), .D(_0626_), .Q(round_key[107]));
    dff _6211_(.RN(_0238_), .SN(1'b1), .CK(clk), .D(_0627_), .Q(round_key[108]));
    dff _6212_(.RN(_0239_), .SN(1'b1), .CK(clk), .D(_0628_), .Q(round_key[109]));
    dff _6213_(.RN(_0240_), .SN(1'b1), .CK(clk), .D(_0629_), .Q(round_key[110]));
    dff _6214_(.RN(_0241_), .SN(1'b1), .CK(clk), .D(_0630_), .Q(round_key[111]));
    dff _6215_(.RN(_0242_), .SN(1'b1), .CK(clk), .D(_0631_), .Q(round_key[112]));
    dff _6216_(.RN(_0243_), .SN(1'b1), .CK(clk), .D(_0632_), .Q(round_key[113]));
    dff _6217_(.RN(_0244_), .SN(1'b1), .CK(clk), .D(_0633_), .Q(round_key[114]));
    dff _6218_(.RN(_0245_), .SN(1'b1), .CK(clk), .D(_0634_), .Q(round_key[115]));
    dff _6219_(.RN(_0246_), .SN(1'b1), .CK(clk), .D(_0635_), .Q(round_key[116]));
    dff _6220_(.RN(_0247_), .SN(1'b1), .CK(clk), .D(_0636_), .Q(round_key[117]));
    dff _6221_(.RN(_0248_), .SN(1'b1), .CK(clk), .D(_0637_), .Q(round_key[118]));
    dff _6222_(.RN(_0249_), .SN(1'b1), .CK(clk), .D(_0638_), .Q(round_key[119]));
    dff _6223_(.RN(_0250_), .SN(1'b1), .CK(clk), .D(_0639_), .Q(round_key[120]));
    dff _6224_(.RN(_0251_), .SN(1'b1), .CK(clk), .D(_0640_), .Q(round_key[121]));
    dff _6225_(.RN(_0252_), .SN(1'b1), .CK(clk), .D(_0641_), .Q(round_key[122]));
    dff _6226_(.RN(_0253_), .SN(1'b1), .CK(clk), .D(_0642_), .Q(round_key[123]));
    dff _6227_(.RN(_0254_), .SN(1'b1), .CK(clk), .D(_0643_), .Q(round_key[124]));
    dff _6228_(.RN(_0255_), .SN(1'b1), .CK(clk), .D(_0644_), .Q(round_key[125]));
    dff _6229_(.RN(_0256_), .SN(1'b1), .CK(clk), .D(_0645_), .Q(round_key[126]));
    dff _6230_(.RN(_0257_), .SN(1'b1), .CK(clk), .D(_0646_), .Q(round_key[127]));
    dff _6231_(.RN(_0258_), .SN(1'b1), .CK(clk), .D(_0647_), .Q(round_counter[0]));
    dff _6232_(.RN(_0259_), .SN(1'b1), .CK(clk), .D(_0648_), .Q(round_counter[1]));
    dff _6233_(.RN(_0260_), .SN(1'b1), .CK(clk), .D(_0649_), .Q(round_counter[2]));
    dff _6234_(.RN(_0261_), .SN(1'b1), .CK(clk), .D(_0650_), .Q(ciphertext[0]));
    dff _6235_(.RN(_0262_), .SN(1'b1), .CK(clk), .D(_0651_), .Q(ciphertext[1]));
    dff _6236_(.RN(_0263_), .SN(1'b1), .CK(clk), .D(_0000_), .Q(encrypting));
    dff _6237_(.RN(_0264_), .SN(1'b1), .CK(clk), .D(_0652_), .Q(ciphertext[2]));
    dff _6238_(.RN(_0265_), .SN(1'b1), .CK(clk), .D(_0653_), .Q(ciphertext[3]));
    dff _6239_(.RN(_0266_), .SN(1'b1), .CK(clk), .D(_0654_), .Q(ciphertext[4]));
    dff _6240_(.RN(_0267_), .SN(1'b1), .CK(clk), .D(_0655_), .Q(ciphertext[5]));
    dff _6241_(.RN(_0268_), .SN(1'b1), .CK(clk), .D(_0656_), .Q(ciphertext[6]));
    dff _6242_(.RN(_0269_), .SN(1'b1), .CK(clk), .D(_0657_), .Q(ciphertext[7]));
    dff _6243_(.RN(_0270_), .SN(1'b1), .CK(clk), .D(_0658_), .Q(ciphertext[8]));
    dff _6244_(.RN(_0271_), .SN(1'b1), .CK(clk), .D(_0659_), .Q(ciphertext[9]));
    dff _6245_(.RN(_0272_), .SN(1'b1), .CK(clk), .D(_0660_), .Q(ciphertext[10]));
    dff _6246_(.RN(_0273_), .SN(1'b1), .CK(clk), .D(_0661_), .Q(ciphertext[11]));
    dff _6247_(.RN(_0274_), .SN(1'b1), .CK(clk), .D(_0662_), .Q(ciphertext[12]));
    dff _6248_(.RN(_0275_), .SN(1'b1), .CK(clk), .D(_0663_), .Q(ciphertext[13]));
    dff _6249_(.RN(_0276_), .SN(1'b1), .CK(clk), .D(_0664_), .Q(ciphertext[14]));
    dff _6250_(.RN(_0277_), .SN(1'b1), .CK(clk), .D(_0665_), .Q(ciphertext[15]));
    dff _6251_(.RN(_0278_), .SN(1'b1), .CK(clk), .D(_0666_), .Q(ciphertext[16]));
    dff _6252_(.RN(_0279_), .SN(1'b1), .CK(clk), .D(_0667_), .Q(ciphertext[17]));
    dff _6253_(.RN(_0280_), .SN(1'b1), .CK(clk), .D(_0668_), .Q(ciphertext[18]));
    dff _6254_(.RN(_0281_), .SN(1'b1), .CK(clk), .D(_0669_), .Q(ciphertext[19]));
    dff _6255_(.RN(_0282_), .SN(1'b1), .CK(clk), .D(_0670_), .Q(ciphertext[20]));
    dff _6256_(.RN(_0283_), .SN(1'b1), .CK(clk), .D(_0671_), .Q(ciphertext[21]));
    dff _6257_(.RN(_0284_), .SN(1'b1), .CK(clk), .D(_0672_), .Q(ciphertext[22]));
    dff _6258_(.RN(_0285_), .SN(1'b1), .CK(clk), .D(_0673_), .Q(ciphertext[23]));
    dff _6259_(.RN(_0286_), .SN(1'b1), .CK(clk), .D(_0674_), .Q(ciphertext[24]));
    dff _6260_(.RN(_0287_), .SN(1'b1), .CK(clk), .D(_0675_), .Q(ciphertext[25]));
    dff _6261_(.RN(_0288_), .SN(1'b1), .CK(clk), .D(_0676_), .Q(ciphertext[26]));
    dff _6262_(.RN(_0289_), .SN(1'b1), .CK(clk), .D(_0677_), .Q(ciphertext[27]));
    dff _6263_(.RN(_0290_), .SN(1'b1), .CK(clk), .D(_0678_), .Q(ciphertext[28]));
    dff _6264_(.RN(_0291_), .SN(1'b1), .CK(clk), .D(_0679_), .Q(ciphertext[29]));
    dff _6265_(.RN(_0292_), .SN(1'b1), .CK(clk), .D(_0680_), .Q(ciphertext[30]));
    dff _6266_(.RN(_0293_), .SN(1'b1), .CK(clk), .D(_0681_), .Q(ciphertext[31]));
    dff _6267_(.RN(_0294_), .SN(1'b1), .CK(clk), .D(_0682_), .Q(ciphertext[32]));
    dff _6268_(.RN(_0295_), .SN(1'b1), .CK(clk), .D(_0683_), .Q(ciphertext[33]));
    dff _6269_(.RN(_0296_), .SN(1'b1), .CK(clk), .D(_0684_), .Q(ciphertext[34]));
    dff _6270_(.RN(_0297_), .SN(1'b1), .CK(clk), .D(_0685_), .Q(ciphertext[35]));
    dff _6271_(.RN(_0298_), .SN(1'b1), .CK(clk), .D(_0686_), .Q(ciphertext[36]));
    dff _6272_(.RN(_0299_), .SN(1'b1), .CK(clk), .D(_0687_), .Q(ciphertext[37]));
    dff _6273_(.RN(_0300_), .SN(1'b1), .CK(clk), .D(_0688_), .Q(ciphertext[38]));
    dff _6274_(.RN(_0301_), .SN(1'b1), .CK(clk), .D(_0689_), .Q(ciphertext[39]));
    dff _6275_(.RN(_0302_), .SN(1'b1), .CK(clk), .D(_0690_), .Q(ciphertext[40]));
    dff _6276_(.RN(_0303_), .SN(1'b1), .CK(clk), .D(_0691_), .Q(ciphertext[41]));
    dff _6277_(.RN(_0304_), .SN(1'b1), .CK(clk), .D(_0692_), .Q(ciphertext[42]));
    dff _6278_(.RN(_0305_), .SN(1'b1), .CK(clk), .D(_0693_), .Q(ciphertext[43]));
    dff _6279_(.RN(_0306_), .SN(1'b1), .CK(clk), .D(_0694_), .Q(ciphertext[44]));
    dff _6280_(.RN(_0307_), .SN(1'b1), .CK(clk), .D(_0695_), .Q(ciphertext[45]));
    dff _6281_(.RN(_0308_), .SN(1'b1), .CK(clk), .D(_0696_), .Q(ciphertext[46]));
    dff _6282_(.RN(_0309_), .SN(1'b1), .CK(clk), .D(_0697_), .Q(ciphertext[47]));
    dff _6283_(.RN(_0310_), .SN(1'b1), .CK(clk), .D(_0698_), .Q(ciphertext[48]));
    dff _6284_(.RN(_0311_), .SN(1'b1), .CK(clk), .D(_0699_), .Q(ciphertext[49]));
    dff _6285_(.RN(_0312_), .SN(1'b1), .CK(clk), .D(_0700_), .Q(ciphertext[50]));
    dff _6286_(.RN(_0313_), .SN(1'b1), .CK(clk), .D(_0701_), .Q(ciphertext[51]));
    dff _6287_(.RN(_0314_), .SN(1'b1), .CK(clk), .D(_0702_), .Q(ciphertext[52]));
    dff _6288_(.RN(_0315_), .SN(1'b1), .CK(clk), .D(_0703_), .Q(ciphertext[53]));
    dff _6289_(.RN(_0316_), .SN(1'b1), .CK(clk), .D(_0704_), .Q(ciphertext[54]));
    dff _6290_(.RN(_0317_), .SN(1'b1), .CK(clk), .D(_0705_), .Q(ciphertext[55]));
    dff _6291_(.RN(_0318_), .SN(1'b1), .CK(clk), .D(_0706_), .Q(ciphertext[56]));
    dff _6292_(.RN(_0319_), .SN(1'b1), .CK(clk), .D(_0707_), .Q(ciphertext[57]));
    dff _6293_(.RN(_0320_), .SN(1'b1), .CK(clk), .D(_0708_), .Q(ciphertext[58]));
    dff _6294_(.RN(_0321_), .SN(1'b1), .CK(clk), .D(_0709_), .Q(ciphertext[59]));
    dff _6295_(.RN(_0322_), .SN(1'b1), .CK(clk), .D(_0710_), .Q(ciphertext[60]));
    dff _6296_(.RN(_0323_), .SN(1'b1), .CK(clk), .D(_0711_), .Q(ciphertext[61]));
    dff _6297_(.RN(_0324_), .SN(1'b1), .CK(clk), .D(_0712_), .Q(ciphertext[62]));
    dff _6298_(.RN(_0325_), .SN(1'b1), .CK(clk), .D(_0713_), .Q(ciphertext[63]));
    dff _6299_(.RN(_0326_), .SN(1'b1), .CK(clk), .D(_0714_), .Q(ciphertext[64]));
    dff _6300_(.RN(_0327_), .SN(1'b1), .CK(clk), .D(_0715_), .Q(ciphertext[65]));
    dff _6301_(.RN(_0328_), .SN(1'b1), .CK(clk), .D(_0716_), .Q(ciphertext[66]));
    dff _6302_(.RN(_0329_), .SN(1'b1), .CK(clk), .D(_0717_), .Q(ciphertext[67]));
    dff _6303_(.RN(_0330_), .SN(1'b1), .CK(clk), .D(_0718_), .Q(ciphertext[68]));
    dff _6304_(.RN(_0331_), .SN(1'b1), .CK(clk), .D(_0719_), .Q(ciphertext[69]));
    dff _6305_(.RN(_0332_), .SN(1'b1), .CK(clk), .D(_0720_), .Q(ciphertext[70]));
    dff _6306_(.RN(_0333_), .SN(1'b1), .CK(clk), .D(_0721_), .Q(ciphertext[71]));
    dff _6307_(.RN(_0334_), .SN(1'b1), .CK(clk), .D(_0722_), .Q(ciphertext[72]));
    dff _6308_(.RN(_0335_), .SN(1'b1), .CK(clk), .D(_0723_), .Q(ciphertext[73]));
    dff _6309_(.RN(_0336_), .SN(1'b1), .CK(clk), .D(_0724_), .Q(ciphertext[74]));
    dff _6310_(.RN(_0337_), .SN(1'b1), .CK(clk), .D(_0725_), .Q(ciphertext[75]));
    dff _6311_(.RN(_0338_), .SN(1'b1), .CK(clk), .D(_0726_), .Q(ciphertext[76]));
    dff _6312_(.RN(_0339_), .SN(1'b1), .CK(clk), .D(_0727_), .Q(ciphertext[77]));
    dff _6313_(.RN(_0340_), .SN(1'b1), .CK(clk), .D(_0728_), .Q(ciphertext[78]));
    dff _6314_(.RN(_0341_), .SN(1'b1), .CK(clk), .D(_0729_), .Q(ciphertext[79]));
    dff _6315_(.RN(_0342_), .SN(1'b1), .CK(clk), .D(_0730_), .Q(ciphertext[80]));
    dff _6316_(.RN(_0343_), .SN(1'b1), .CK(clk), .D(_0731_), .Q(ciphertext[81]));
    dff _6317_(.RN(_0344_), .SN(1'b1), .CK(clk), .D(_0732_), .Q(ciphertext[82]));
    dff _6318_(.RN(_0345_), .SN(1'b1), .CK(clk), .D(_0733_), .Q(ciphertext[83]));
    dff _6319_(.RN(_0346_), .SN(1'b1), .CK(clk), .D(_0734_), .Q(ciphertext[84]));
    dff _6320_(.RN(_0347_), .SN(1'b1), .CK(clk), .D(_0735_), .Q(ciphertext[85]));
    dff _6321_(.RN(_0348_), .SN(1'b1), .CK(clk), .D(_0736_), .Q(ciphertext[86]));
    dff _6322_(.RN(_0349_), .SN(1'b1), .CK(clk), .D(_0737_), .Q(ciphertext[87]));
    dff _6323_(.RN(_0350_), .SN(1'b1), .CK(clk), .D(_0738_), .Q(ciphertext[88]));
    dff _6324_(.RN(_0351_), .SN(1'b1), .CK(clk), .D(_0739_), .Q(ciphertext[89]));
    dff _6325_(.RN(_0352_), .SN(1'b1), .CK(clk), .D(_0740_), .Q(ciphertext[90]));
    dff _6326_(.RN(_0353_), .SN(1'b1), .CK(clk), .D(_0741_), .Q(ciphertext[91]));
    dff _6327_(.RN(_0354_), .SN(1'b1), .CK(clk), .D(_0742_), .Q(ciphertext[92]));
    dff _6328_(.RN(_0355_), .SN(1'b1), .CK(clk), .D(_0743_), .Q(ciphertext[93]));
    dff _6329_(.RN(_0356_), .SN(1'b1), .CK(clk), .D(_0744_), .Q(ciphertext[94]));
    dff _6330_(.RN(_0357_), .SN(1'b1), .CK(clk), .D(_0745_), .Q(ciphertext[95]));
    dff _6331_(.RN(_0358_), .SN(1'b1), .CK(clk), .D(_0746_), .Q(ciphertext[96]));
    dff _6332_(.RN(_0359_), .SN(1'b1), .CK(clk), .D(_0747_), .Q(ciphertext[97]));
    dff _6333_(.RN(_0360_), .SN(1'b1), .CK(clk), .D(_0748_), .Q(ciphertext[98]));
    dff _6334_(.RN(_0361_), .SN(1'b1), .CK(clk), .D(_0749_), .Q(ciphertext[99]));
    dff _6335_(.RN(_0362_), .SN(1'b1), .CK(clk), .D(_0750_), .Q(ciphertext[100]));
    dff _6336_(.RN(_0363_), .SN(1'b1), .CK(clk), .D(_0751_), .Q(ciphertext[101]));
    dff _6337_(.RN(_0364_), .SN(1'b1), .CK(clk), .D(_0752_), .Q(ciphertext[102]));
    dff _6338_(.RN(_0365_), .SN(1'b1), .CK(clk), .D(_0753_), .Q(ciphertext[103]));
    dff _6339_(.RN(_0366_), .SN(1'b1), .CK(clk), .D(_0754_), .Q(ciphertext[104]));
    dff _6340_(.RN(_0367_), .SN(1'b1), .CK(clk), .D(_0755_), .Q(ciphertext[105]));
    dff _6341_(.RN(_0368_), .SN(1'b1), .CK(clk), .D(_0756_), .Q(ciphertext[106]));
    dff _6342_(.RN(_0369_), .SN(1'b1), .CK(clk), .D(_0757_), .Q(ciphertext[107]));
    dff _6343_(.RN(_0370_), .SN(1'b1), .CK(clk), .D(_0758_), .Q(ciphertext[108]));
    dff _6344_(.RN(_0371_), .SN(1'b1), .CK(clk), .D(_0759_), .Q(ciphertext[109]));
    dff _6345_(.RN(_0372_), .SN(1'b1), .CK(clk), .D(_0760_), .Q(ciphertext[110]));
    dff _6346_(.RN(_0373_), .SN(1'b1), .CK(clk), .D(_0761_), .Q(ciphertext[111]));
    dff _6347_(.RN(_0374_), .SN(1'b1), .CK(clk), .D(_0762_), .Q(ciphertext[112]));
    dff _6348_(.RN(_0375_), .SN(1'b1), .CK(clk), .D(_0763_), .Q(ciphertext[113]));
    dff _6349_(.RN(_0376_), .SN(1'b1), .CK(clk), .D(_0764_), .Q(ciphertext[114]));
    dff _6350_(.RN(_0377_), .SN(1'b1), .CK(clk), .D(_0765_), .Q(ciphertext[115]));
    dff _6351_(.RN(_0378_), .SN(1'b1), .CK(clk), .D(_0766_), .Q(ciphertext[116]));
    dff _6352_(.RN(_0379_), .SN(1'b1), .CK(clk), .D(_0767_), .Q(ciphertext[117]));
    dff _6353_(.RN(_0380_), .SN(1'b1), .CK(clk), .D(_0768_), .Q(ciphertext[118]));
    dff _6354_(.RN(_0381_), .SN(1'b1), .CK(clk), .D(_0769_), .Q(ciphertext[119]));
    dff _6355_(.RN(_0382_), .SN(1'b1), .CK(clk), .D(_0770_), .Q(ciphertext[120]));
    dff _6356_(.RN(_0383_), .SN(1'b1), .CK(clk), .D(_0771_), .Q(ciphertext[121]));
    dff _6357_(.RN(_0384_), .SN(1'b1), .CK(clk), .D(_0772_), .Q(ciphertext[122]));
    dff _6358_(.RN(_0385_), .SN(1'b1), .CK(clk), .D(_0773_), .Q(ciphertext[123]));
    dff _6359_(.RN(_0386_), .SN(1'b1), .CK(clk), .D(_0774_), .Q(ciphertext[124]));
    dff _6360_(.RN(_0387_), .SN(1'b1), .CK(clk), .D(_0775_), .Q(ciphertext[125]));
    dff _6361_(.RN(_0388_), .SN(1'b1), .CK(clk), .D(_0776_), .Q(ciphertext[126]));
    dff _6362_(.RN(_0389_), .SN(1'b1), .CK(clk), .D(_0777_), .Q(ciphertext[127]));
endmodule