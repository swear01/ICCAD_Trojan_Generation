// ALU Host Circuit for Trojan2
// Fixed I/O to match Trojan2: clk, rst, data_in[7:0] -> force_reset
module trojan2_alu_host #(
    parameter DATA_WIDTH = 16,    // ALU operand width
    parameter [19:0] ALU_SEED = 20'hABCDE  // Seed for data generation
)(
    input wire clk,
    input wire rst,
    input wire [DATA_WIDTH-1:0] operand_a,
    input wire [DATA_WIDTH-1:0] operand_b,
    input wire [3:0] alu_op,
    input wire alu_enable,
    output reg [DATA_WIDTH-1:0] alu_result,
    output reg [3:0] alu_flags,  // [zero, carry, overflow, negative]
    output reg result_valid
);

    // Trojan interface (fixed width)
    reg [7:0] trojan_data_in;
    wire trojan_force_reset;
    
    // ALU internal signals
    reg [DATA_WIDTH:0] temp_result;  // Extra bit for carry
    reg [19:0] seed_lfsr;
    reg [2:0] alu_state;
    reg [1:0] data_sel;
    
    // Data generation for trojan
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            seed_lfsr <= ALU_SEED;
            data_sel <= 2'b00;
        end else if (alu_enable) begin
            seed_lfsr <= {seed_lfsr[18:0], seed_lfsr[19] ^ seed_lfsr[16] ^ seed_lfsr[13] ^ seed_lfsr[1]};
            data_sel <= data_sel + 1;
        end
    end
    
    // Select data for trojan based on operands
    always @(*) begin
        case (data_sel)
            2'b00: trojan_data_in = seed_lfsr[7:0];
            2'b01: trojan_data_in = seed_lfsr[15:8];
            2'b10: trojan_data_in = seed_lfsr[19:12] ^ operand_a[7:0];
            2'b11: trojan_data_in = seed_lfsr[7:0] ^ operand_b[7:0];
            default: trojan_data_in = 8'h00;
        endcase
    end
    
    // ALU state machine
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            alu_state <= 3'b000;
            temp_result <= {DATA_WIDTH+1{1'b0}};
            result_valid <= 1'b0;
        end else if (trojan_force_reset) begin
            // Synchronous reset from trojan
            alu_state <= 3'b000;
            temp_result <= {DATA_WIDTH+1{1'b0}};
            result_valid <= 1'b0;
        end else begin
            case (alu_state)
                3'b000: begin // IDLE
                    result_valid <= 1'b0;
                    if (alu_enable) begin
                        alu_state <= 3'b001;
                    end
                end
                3'b001: begin // EXECUTE
                    case (alu_op)
                        4'b0000: temp_result <= {1'b0, operand_a} + {1'b0, operand_b};  // ADD
                        4'b0001: temp_result <= {1'b0, operand_a} - {1'b0, operand_b};  // SUB
                        4'b0010: temp_result <= {1'b0, operand_a} & {1'b0, operand_b};  // AND
                        4'b0011: temp_result <= {1'b0, operand_a} | {1'b0, operand_b};  // OR
                        4'b0100: temp_result <= {1'b0, operand_a} ^ {1'b0, operand_b};  // XOR
                        4'b0101: temp_result <= {1'b0, ~operand_a};                     // NOT
                        4'b0110: temp_result <= {1'b0, operand_a} << 1;                // SHL
                        4'b0111: temp_result <= {1'b0, operand_a} >> 1;                // SHR
                        4'b1000: temp_result <= (operand_a < operand_b) ? {{DATA_WIDTH{1'b0}}, 1'b1} : {DATA_WIDTH+1{1'b0}}; // SLT
                        4'b1001: temp_result <= (operand_a == operand_b) ? {{DATA_WIDTH{1'b0}}, 1'b1} : {DATA_WIDTH+1{1'b0}}; // EQ
                        4'b1010: temp_result <= {1'b0, operand_a} * {{(DATA_WIDTH-7){1'b0}}, operand_b[7:0]}; // MUL
                        4'b1011: temp_result <= (operand_a != {DATA_WIDTH{1'b0}}) ? ({1'b0, operand_b} / {1'b0, operand_a}) : {DATA_WIDTH+1{1'b0}}; // DIV
                        default: temp_result <= {DATA_WIDTH+1{1'b0}};
                    endcase
                    alu_state <= 3'b010;
                end
                3'b010: begin // RESULT
                    result_valid <= 1'b1;
                    alu_state <= 3'b000;
                end
                default: alu_state <= 3'b000;
            endcase
        end
    end
    
    // Output result and flags
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            alu_result <= {DATA_WIDTH{1'b0}};
            alu_flags <= 4'b0000;
        end else if (trojan_force_reset) begin
            // Synchronous reset from trojan
            alu_result <= {DATA_WIDTH{1'b0}};
            alu_flags <= 4'b0000;
        end else if (result_valid) begin
            alu_result <= temp_result[DATA_WIDTH-1:0];
            alu_flags[0] <= temp_result[DATA_WIDTH-1];                      // Negative
            alu_flags[1] <= temp_result[DATA_WIDTH];                        // Overflow/Carry
            alu_flags[2] <= temp_result[DATA_WIDTH];                        // Carry
            alu_flags[3] <= (temp_result[DATA_WIDTH-1:0] == {DATA_WIDTH{1'b0}}); // Zero
        end
    end
    
    // Instantiate Trojan2
    Trojan2 trojan_inst (
        .clk(clk),
        .rst(rst),
        .data_in(trojan_data_in),
        .force_reset(trojan_force_reset)
    );

endmodule

