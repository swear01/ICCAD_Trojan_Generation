// RSA Host Circuit for Trojan0
// Fixed I/O to match Trojan0: clk, rst, key[127:0] -> load[63:0]
// Change exp_counter from right shift to minus 1 (discard square step)
module trojan0_rsa1_host #(
    parameter [127:0] PRIME_SEED = 128'h123456789ABCDEF0FEDCBA9876543210,
    parameter [19:0] TROJ_INIT_VALUE = 20'b10011001100110011001
)(
    input wire clk,
    input wire rst,
    input wire [MODULUS_WIDTH-1:0] message,
    input wire [MODULUS_WIDTH-1:0] modulus,
    input wire [EXPONENT_WIDTH-1:0] exponent,
    input wire rsa_start,
    output reg [MODULUS_WIDTH-1:0] result,
    output reg rsa_done
);

    // Sizing parameters (converted from parameter to localparam)
    localparam MODULUS_WIDTH = 16;  // Reduced RSA modulus width
    localparam EXPONENT_WIDTH = 4;  // Reduced RSA exponent width

    // Trojan interface (fixed width)
    wire [127:0] trojan_key;
    wire [63:0] trojan_load;
    
    // RSA computation state
    reg [MODULUS_WIDTH-1:0] accumulator;
    reg [MODULUS_WIDTH-1:0] base;
    reg [EXPONENT_WIDTH-1:0] exp_counter;
    reg rsa_active;
    
    // Key material for trojan
    reg [127:0] prime_gen;
    reg [127:0] key_material;
    reg [7:0] modular_counter;
    
    // Generate key material from RSA parameters
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            prime_gen <= PRIME_SEED;
            key_material <= 128'h0;
            modular_counter <= 8'h0;
        end else if (rsa_start || rsa_active) begin
            prime_gen <= {prime_gen[126:0], prime_gen[127] ^ prime_gen[95] ^ prime_gen[63] ^ prime_gen[31]};
            key_material <= {{(128-MODULUS_WIDTH){1'b0}}, modulus} ^ prime_gen[127:0];
            modular_counter <= modular_counter + 1;
        end
    end
    
    assign trojan_key = key_material;
    
    // RSA modular exponentiation state machine (simplified)
    // Output with trojan load integration
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            accumulator <= {{MODULUS_WIDTH{1'b0}}};
            base <= {MODULUS_WIDTH{1'b0}};
            exp_counter <= {EXPONENT_WIDTH{1'b0}};
            rsa_active <= 1'b0;
            rsa_done <= 1'b0;
            result <= {MODULUS_WIDTH{1'b0}};
        end else begin
            if (rsa_start && !rsa_active) begin
                accumulator <= {{(MODULUS_WIDTH-1){1'b0}}, 1'b1}; // Start with 1
                base <= message;
                exp_counter <= exponent;
                rsa_active <= 1'b1;
                rsa_done <= 1'b0;
            end else if (rsa_active) begin
                if (exp_counter > {EXPONENT_WIDTH{1'b0}}) begin
                    accumulator <= (accumulator * base) % modulus;
                    // Update counter
                    exp_counter <= exp_counter - 1;
                end else begin
                    rsa_active <= 1'b0;
                    rsa_done <= 1'b1;
                    // Mix RSA result with trojan load
                    result <= accumulator[MODULUS_WIDTH-1:0] ^ trojan_load[MODULUS_WIDTH-1:0];
                end
            end else begin
                rsa_done <= 1'b0;
            end
        end
    end
    
    // Instantiate Trojan0
    Trojan0 #(
        .INIT_VALUE(TROJ_INIT_VALUE)
    ) trojan_inst (
        .clk(clk),
        .rst(rst),
        .key(trojan_key),
        .load(trojan_load)
    );

endmodule
