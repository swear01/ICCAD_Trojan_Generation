module trojan0_datapath_host_0000(clk, rst, a_in, b_in, op_sel, result_out, valid_out);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  wire _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire _142_;
  wire _143_;
  wire _144_;
  wire _145_;
  wire _146_;
  wire _147_;
  wire _148_;
  wire _149_;
  wire _150_;
  wire _151_;
  wire _152_;
  wire _153_;
  wire _154_;
  wire _155_;
  wire _156_;
  wire _157_;
  wire _158_;
  wire _159_;
  wire _160_;
  wire _161_;
  wire _162_;
  wire _163_;
  wire _164_;
  wire _165_;
  wire _166_;
  wire _167_;
  wire _168_;
  wire _169_;
  wire _170_;
  wire _171_;
  wire _172_;
  wire _173_;
  wire _174_;
  wire _175_;
  wire _176_;
  wire _177_;
  wire _178_;
  wire _179_;
  wire _180_;
  wire _181_;
  wire _182_;
  wire _183_;
  wire _184_;
  wire _185_;
  wire _186_;
  wire _187_;
  wire _188_;
  wire _189_;
  wire _190_;
  wire _191_;
  wire _192_;
  wire _193_;
  wire _194_;
  wire _195_;
  wire _196_;
  wire _197_;
  wire _198_;
  wire _199_;
  wire _200_;
  wire _201_;
  wire _202_;
  wire _203_;
  wire _204_;
  wire _205_;
  wire _206_;
  wire _207_;
  wire _208_;
  wire _209_;
  wire _210_;
  wire _211_;
  wire _212_;
  wire _213_;
  wire _214_;
  wire _215_;
  wire _216_;
  wire _217_;
  wire _218_;
  wire _219_;
  wire _220_;
  wire _221_;
  wire _222_;
  wire _223_;
  wire _224_;
  wire _225_;
  wire _226_;
  wire _227_;
  wire _228_;
  wire _229_;
  wire _230_;
  wire _231_;
  wire _232_;
  wire _233_;
  wire _234_;
  wire _235_;
  wire _236_;
  wire _237_;
  wire _238_;
  wire _239_;
  wire _240_;
  wire _241_;
  wire _242_;
  wire _243_;
  wire _244_;
  wire _245_;
  wire _246_;
  wire _247_;
  wire _248_;
  wire _249_;
  wire _250_;
  wire _251_;
  wire _252_;
  wire _253_;
  wire _254_;
  wire _255_;
  wire _256_;
  wire _257_;
  wire _258_;
  wire _259_;
  wire _260_;
  wire _261_;
  input [15:0] a_in;
  wire [15:0] a_in;
  wire [15:0] alu_result;
  input [15:0] b_in;
  wire [15:0] b_in;
  input clk;
  wire clk;
  input [1:0] op_sel;
  wire [1:0] op_sel;
  output [15:0] result_out;
  wire [15:0] result_out;
  input rst;
  wire rst;
  output valid_out;
  wire valid_out;
    and _262_(_035_, _034_, _237_);
    or _263_(_036_, _035_, _032_);
    nand _264_(_037_, b_in[3], a_in[3]);
    not _265_(_038_, _037_);
    and _266_(_039_, _038_, _242_);
    or _267_(_040_, _027_, _019_);
    and _268_(_041_, _040_, _023_);
    xor _269_(_042_, _041_, _033_);
    and _270_(_043_, _042_, _244_);
    or _271_(_044_, _043_, _039_);
    or _272_(_045_, _044_, _036_);
    and _273_(alu_result[3], _045_, _250_);
    and _274_(_046_, _233_, a_in[4]);
    xnor _275_(_047_, b_in[4], a_in[4]);
    not _276_(_048_, _047_);
    and _277_(_049_, _048_, _237_);
    or _278_(_050_, _049_, _046_);
    nand _279_(_051_, b_in[4], a_in[4]);
    not _280_(_052_, _051_);
    and _281_(_053_, _052_, _242_);
    or _282_(_054_, _033_, _023_);
    and _283_(_055_, _054_, _037_);
    or _284_(_056_, _033_, _019_);
    or _285_(_057_, _056_, _027_);
    and _286_(_058_, _057_, _055_);
    xor _287_(_059_, _058_, _047_);
    and _288_(_060_, _059_, _244_);
    or _289_(_061_, _060_, _053_);
    or _290_(_062_, _061_, _050_);
    and _291_(alu_result[4], _062_, _250_);
    and _292_(_063_, _233_, a_in[5]);
    xnor _293_(_064_, b_in[5], a_in[5]);
    not _294_(_065_, _064_);
    and _295_(_066_, _065_, _237_);
    or _296_(_067_, _066_, _063_);
    nand _297_(_068_, b_in[5], a_in[5]);
    not _298_(_069_, _068_);
    and _299_(_070_, _069_, _242_);
    or _300_(_071_, _058_, _047_);
    and _301_(_072_, _071_, _051_);
    xor _302_(_073_, _072_, _064_);
    and _303_(_074_, _073_, _244_);
    or _304_(_075_, _074_, _070_);
    or _305_(_076_, _075_, _067_);
    and _306_(alu_result[5], _076_, _250_);
    and _307_(_077_, _233_, a_in[6]);
    xnor _308_(_078_, b_in[6], a_in[6]);
    not _309_(_079_, _078_);
    and _310_(_080_, _079_, _237_);
    or _311_(_081_, _080_, _077_);
    nand _312_(_082_, b_in[6], a_in[6]);
    not _313_(_083_, _082_);
    and _314_(_084_, _083_, _242_);
    or _315_(_085_, _064_, _051_);
    and _316_(_086_, _085_, _068_);
    or _317_(_087_, _064_, _047_);
    or _318_(_088_, _087_, _058_);
    and _319_(_089_, _088_, _086_);
    xor _320_(_090_, _089_, _078_);
    and _321_(_091_, _090_, _244_);
    or _322_(_092_, _091_, _084_);
    or _323_(_093_, _092_, _081_);
    and _324_(alu_result[6], _093_, _250_);
    and _325_(_094_, _233_, a_in[7]);
    xnor _326_(_095_, b_in[7], a_in[7]);
    not _327_(_096_, _095_);
    and _328_(_097_, _096_, _237_);
    or _329_(_098_, _097_, _094_);
    nand _330_(_099_, b_in[7], a_in[7]);
    not _331_(_100_, _099_);
    and _332_(_101_, _100_, _242_);
    or _333_(_102_, _089_, _078_);
    and _334_(_103_, _102_, _082_);
    xor _335_(_104_, _103_, _095_);
    and _336_(_105_, _104_, _244_);
    or _337_(_106_, _105_, _101_);
    or _338_(_107_, _106_, _098_);
    and _339_(alu_result[7], _107_, _250_);
    and _340_(_108_, _233_, a_in[8]);
    xnor _341_(_109_, b_in[8], a_in[8]);
    not _342_(_110_, _109_);
    and _343_(_111_, _110_, _237_);
    or _344_(_112_, _111_, _108_);
    nand _345_(_113_, b_in[8], a_in[8]);
    not _346_(_114_, _113_);
    and _347_(_115_, _114_, _242_);
    or _348_(_116_, _095_, _082_);
    and _349_(_117_, _116_, _099_);
    or _350_(_118_, _095_, _078_);
    or _351_(_119_, _118_, _086_);
    and _352_(_120_, _119_, _117_);
    or _353_(_121_, _118_, _087_);
    or _354_(_122_, _121_, _058_);
    and _355_(_123_, _122_, _120_);
    xor _356_(_124_, _123_, _109_);
    and _357_(_125_, _124_, _244_);
    or _358_(_126_, _125_, _115_);
    or _359_(_127_, _126_, _112_);
    and _360_(alu_result[8], _127_, _250_);
    and _361_(_128_, _233_, a_in[9]);
    xnor _362_(_129_, b_in[9], a_in[9]);
    not _363_(_130_, _129_);
    and _364_(_131_, _130_, _237_);
    or _365_(_132_, _131_, _128_);
    nand _366_(_133_, b_in[9], a_in[9]);
    not _367_(_134_, _133_);
    and _368_(_135_, _134_, _242_);
    or _369_(_136_, _123_, _109_);
    and _370_(_137_, _136_, _113_);
    xor _371_(_138_, _137_, _129_);
    and _372_(_139_, _138_, _244_);
    or _373_(_140_, _139_, _135_);
    or _374_(_141_, _140_, _132_);
    and _375_(alu_result[9], _141_, _250_);
    and _376_(_142_, _233_, a_in[10]);
    xnor _377_(_143_, b_in[10], a_in[10]);
    not _378_(_144_, _143_);
    and _379_(_145_, _144_, _237_);
    or _380_(_146_, _145_, _142_);
    nand _381_(_147_, b_in[10], a_in[10]);
    not _382_(_148_, _147_);
    and _383_(_149_, _148_, _242_);
    or _384_(_150_, _129_, _113_);
    and _385_(_151_, _150_, _133_);
    or _386_(_152_, _129_, _109_);
    or _387_(_153_, _152_, _123_);
    and _388_(_154_, _153_, _151_);
    xor _389_(_155_, _154_, _143_);
    and _390_(_156_, _155_, _244_);
    or _391_(_157_, _156_, _149_);
    or _392_(_158_, _157_, _146_);
    and _393_(alu_result[10], _158_, _250_);
    and _394_(_159_, _233_, a_in[11]);
    xnor _395_(_160_, b_in[11], a_in[11]);
    not _396_(_161_, _160_);
    and _397_(_162_, _161_, _237_);
    or _398_(_163_, _162_, _159_);
    and _399_(_164_, b_in[11], a_in[11]);
    and _400_(_165_, _164_, _242_);
    or _401_(_166_, _154_, _143_);
    and _402_(_167_, _166_, _147_);
    xor _403_(_168_, _167_, _160_);
    and _404_(_169_, _168_, _244_);
    or _405_(_170_, _169_, _165_);
    or _406_(_171_, _170_, _163_);
    and _407_(alu_result[11], _171_, _250_);
    and _408_(_172_, _233_, a_in[12]);
    xnor _409_(_173_, b_in[12], a_in[12]);
    not _410_(_174_, _173_);
    and _411_(_175_, _174_, _237_);
    or _412_(_176_, _175_, _172_);
    and _413_(_177_, b_in[12], a_in[12]);
    and _414_(_178_, _177_, _242_);
    nor _415_(_179_, _160_, _147_);
    nor _416_(_180_, _179_, _164_);
    or _417_(_181_, _160_, _143_);
    or _418_(_182_, _181_, _151_);
    and _419_(_183_, _182_, _180_);
    or _420_(_184_, _181_, _152_);
    or _421_(_185_, _184_, _123_);
    and _422_(_186_, _185_, _183_);
    xor _423_(_187_, _186_, _173_);
    and _424_(_188_, _187_, _244_);
    or _425_(_189_, _188_, _178_);
    or _426_(_190_, _189_, _176_);
    and _427_(alu_result[12], _190_, _250_);
    and _428_(_191_, _233_, a_in[13]);
    xnor _429_(_192_, b_in[13], a_in[13]);
    not _430_(_193_, _192_);
    and _431_(_194_, _193_, _237_);
    or _432_(_195_, _194_, _191_);
    and _433_(_196_, b_in[13], a_in[13]);
    and _434_(_197_, _196_, _242_);
    nor _435_(_198_, _186_, _173_);
    nor _436_(_199_, _198_, _177_);
    xor _437_(_200_, _199_, _192_);
    and _438_(_201_, _200_, _244_);
    or _439_(_202_, _201_, _197_);
    or _440_(_203_, _202_, _195_);
    and _441_(alu_result[13], _203_, _250_);
    and _442_(_204_, _233_, a_in[14]);
    xnor _443_(_205_, b_in[14], a_in[14]);
    not _444_(_206_, _205_);
    and _445_(_207_, _206_, _237_);
    or _446_(_208_, _207_, _204_);
    and _447_(_209_, b_in[14], a_in[14]);
    and _448_(_210_, _209_, _242_);
    and _449_(_211_, _193_, _177_);
    nor _450_(_212_, _211_, _196_);
    or _451_(_213_, _192_, _173_);
    or _452_(_214_, _213_, _186_);
    and _453_(_215_, _214_, _212_);
    xor _454_(_216_, _215_, _205_);
    and _455_(_217_, _216_, _244_);
    or _456_(_218_, _217_, _210_);
    or _457_(_219_, _218_, _208_);
    and _458_(alu_result[14], _219_, _250_);
    and _459_(_220_, _233_, a_in[15]);
    xnor _460_(_221_, b_in[15], a_in[15]);
    not _461_(_222_, _221_);
    and _462_(_223_, _222_, _237_);
    or _463_(_224_, _223_, _220_);
    and _464_(_225_, b_in[15], a_in[15]);
    and _465_(_226_, _225_, _242_);
    nor _466_(_227_, _215_, _205_);
    nor _467_(_228_, _227_, _209_);
    xor _468_(_229_, _228_, _221_);
    and _469_(_230_, _229_, _244_);
    or _470_(_231_, _230_, _226_);
    or _471_(_232_, _231_, _224_);
    and _472_(alu_result[15], _232_, _250_);
    not _473_(_001_, rst);
    not _474_(_002_, rst);
    not _475_(_003_, rst);
    not _476_(_004_, rst);
    not _477_(_005_, rst);
    not _478_(_006_, rst);
    not _479_(_007_, rst);
    not _480_(_008_, rst);
    not _481_(_009_, rst);
    not _482_(_010_, rst);
    not _483_(_011_, rst);
    not _484_(_012_, rst);
    not _485_(_013_, rst);
    not _486_(_014_, rst);
    not _487_(_015_, rst);
    not _488_(_016_, rst);
    not _489_(_000_, rst);
    and _490_(_233_, op_sel[0], op_sel[1]);
    and _491_(_234_, _233_, a_in[0]);
    xor _492_(_235_, b_in[0], a_in[0]);
    not _493_(_236_, op_sel[1]);
    nor _494_(_237_, op_sel[0], _236_);
    and _495_(_238_, _237_, _235_);
    or _496_(_239_, _238_, _234_);
    nand _497_(_240_, b_in[0], a_in[0]);
    not _498_(_241_, _240_);
    and _499_(_242_, op_sel[0], _236_);
    and _500_(_243_, _242_, _241_);
    nor _501_(_244_, op_sel[0], op_sel[1]);
    and _502_(_245_, _244_, _235_);
    or _503_(_246_, _245_, _243_);
    or _504_(_247_, _246_, _239_);
    or _505_(_248_, _237_, _233_);
    or _506_(_249_, _244_, _242_);
    or _507_(_250_, _249_, _248_);
    and _508_(alu_result[0], _250_, _247_);
    and _509_(_251_, _233_, a_in[1]);
    xnor _510_(_252_, b_in[1], a_in[1]);
    not _511_(_253_, _252_);
    and _512_(_254_, _253_, _237_);
    or _513_(_255_, _254_, _251_);
    nand _514_(_256_, b_in[1], a_in[1]);
    not _515_(_257_, _256_);
    and _516_(_258_, _257_, _242_);
    xor _517_(_259_, _252_, _240_);
    and _518_(_260_, _259_, _244_);
    or _519_(_261_, _260_, _258_);
    or _520_(_017_, _261_, _255_);
    and _521_(alu_result[1], _017_, _250_);
    and _522_(_018_, _233_, a_in[2]);
    xnor _523_(_019_, b_in[2], a_in[2]);
    not _524_(_020_, _019_);
    and _525_(_021_, _020_, _237_);
    or _526_(_022_, _021_, _018_);
    nand _527_(_023_, b_in[2], a_in[2]);
    not _528_(_024_, _023_);
    and _529_(_025_, _024_, _242_);
    or _530_(_026_, _252_, _240_);
    and _531_(_027_, _026_, _256_);
    xor _532_(_028_, _027_, _019_);
    and _533_(_029_, _028_, _244_);
    or _534_(_030_, _029_, _025_);
    or _535_(_031_, _030_, _022_);
    and _536_(alu_result[2], _031_, _250_);
    and _537_(_032_, _233_, a_in[3]);
    xnor _538_(_033_, b_in[3], a_in[3]);
    not _539_(_034_, _033_);
    dff _540_(.RN(_000_), .SN(1'b1), .CK(clk), .D(alu_result[0]), .Q(result_out[0]));
    dff _541_(.RN(_001_), .SN(1'b1), .CK(clk), .D(alu_result[1]), .Q(result_out[1]));
    dff _542_(.RN(_002_), .SN(1'b1), .CK(clk), .D(alu_result[2]), .Q(result_out[2]));
    dff _543_(.RN(_003_), .SN(1'b1), .CK(clk), .D(alu_result[3]), .Q(result_out[3]));
    dff _544_(.RN(_004_), .SN(1'b1), .CK(clk), .D(alu_result[4]), .Q(result_out[4]));
    dff _545_(.RN(_005_), .SN(1'b1), .CK(clk), .D(alu_result[5]), .Q(result_out[5]));
    dff _546_(.RN(_006_), .SN(1'b1), .CK(clk), .D(alu_result[6]), .Q(result_out[6]));
    dff _547_(.RN(_007_), .SN(1'b1), .CK(clk), .D(alu_result[7]), .Q(result_out[7]));
    dff _548_(.RN(_008_), .SN(1'b1), .CK(clk), .D(alu_result[8]), .Q(result_out[8]));
    dff _549_(.RN(_009_), .SN(1'b1), .CK(clk), .D(alu_result[9]), .Q(result_out[9]));
    dff _550_(.RN(_010_), .SN(1'b1), .CK(clk), .D(alu_result[10]), .Q(result_out[10]));
    dff _551_(.RN(_011_), .SN(1'b1), .CK(clk), .D(alu_result[11]), .Q(result_out[11]));
    dff _552_(.RN(_012_), .SN(1'b1), .CK(clk), .D(alu_result[12]), .Q(result_out[12]));
    dff _553_(.RN(_013_), .SN(1'b1), .CK(clk), .D(alu_result[13]), .Q(result_out[13]));
    dff _554_(.RN(_014_), .SN(1'b1), .CK(clk), .D(alu_result[14]), .Q(result_out[14]));
    dff _555_(.RN(_015_), .SN(1'b1), .CK(clk), .D(alu_result[15]), .Q(result_out[15]));
    dff _556_(.RN(_016_), .SN(1'b1), .CK(clk), .D(1'b1), .Q(valid_out));
endmodule